module plru_decoder (
	way_idx,
	lru_data,
	lru_mask
);
	// Trace: src/VX_cache_repl.sv:2:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_repl.sv:3:15
	parameter WAY_IDX_BITS = $clog2(NUM_WAYS);
	// Trace: src/VX_cache_repl.sv:4:15
	parameter WAY_IDX_WIDTH = (WAY_IDX_BITS > 0 ? WAY_IDX_BITS : 1);
	// Trace: src/VX_cache_repl.sv:6:5
	input wire [WAY_IDX_WIDTH - 1:0] way_idx;
	// Trace: src/VX_cache_repl.sv:7:5
	output wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] lru_data;
	// Trace: src/VX_cache_repl.sv:8:5
	output wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] lru_mask;
	// Trace: src/VX_cache_repl.sv:10:5
	generate
		if (NUM_WAYS > 1) begin : g_dec
			// Trace: src/VX_cache_repl.sv:11:9
			wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] data;
			// Trace: src/VX_cache_repl.sv:12:9
			wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] mask;
			genvar _gv_i_1;
			for (_gv_i_1 = 0; _gv_i_1 < (NUM_WAYS - 1); _gv_i_1 = _gv_i_1 + 1) begin : g_i
				localparam i = _gv_i_1;
				if (i == 0) begin : g_i_0
					// Trace: src/VX_cache_repl.sv:15:17
					assign mask[i] = 1'b1;
				end
				else if ((i % 2) == 1) begin : g_i_odd
					// Trace: src/VX_cache_repl.sv:17:17
					assign mask[i] = mask[(i - 1) / 2] & ~way_idx[(WAY_IDX_BITS - $clog2(i + 2)) + 1];
				end
				else begin : g_i_even
					// Trace: src/VX_cache_repl.sv:19:17
					assign mask[i] = mask[(i - 2) / 2] & way_idx[(WAY_IDX_BITS - $clog2(i + 2)) + 1];
				end
				// Trace: src/VX_cache_repl.sv:21:13
				assign data[i] = ~way_idx[WAY_IDX_BITS - $clog2(i + 2)];
			end
			// Trace: src/VX_cache_repl.sv:23:9
			assign lru_data = data;
			// Trace: src/VX_cache_repl.sv:24:9
			assign lru_mask = mask;
		end
		else begin : g_no_dec
			// Trace: src/VX_cache_repl.sv:26:9
			assign lru_data = 1'sb0;
			// Trace: src/VX_cache_repl.sv:27:9
			assign lru_mask = 1'sb0;
		end
	endgenerate
endmodule
module plru_encoder (
	lru_in,
	way_idx
);
	// Trace: src/VX_cache_repl.sv:31:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_repl.sv:32:15
	parameter WAY_IDX_BITS = $clog2(NUM_WAYS);
	// Trace: src/VX_cache_repl.sv:33:15
	parameter WAY_IDX_WIDTH = (WAY_IDX_BITS > 0 ? WAY_IDX_BITS : 1);
	// Trace: src/VX_cache_repl.sv:35:5
	input wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] lru_in;
	// Trace: src/VX_cache_repl.sv:36:5
	output wire [WAY_IDX_WIDTH - 1:0] way_idx;
	// Trace: src/VX_cache_repl.sv:38:5
	generate
		if (NUM_WAYS > 1) begin : g_enc
			// Trace: src/VX_cache_repl.sv:39:9
			wire [WAY_IDX_BITS - 1:0] tmp;
			genvar _gv_i_2;
			for (_gv_i_2 = 0; _gv_i_2 < WAY_IDX_BITS; _gv_i_2 = _gv_i_2 + 1) begin : g_i
				localparam i = _gv_i_2;
				if (i == 0) begin : g_i_0
					// Trace: src/VX_cache_repl.sv:42:17
					assign tmp[WAY_IDX_WIDTH - 1] = lru_in[0];
				end
				else begin : g_i_n
					// Trace: src/VX_cache_repl.sv:44:17
					VX_mux #(.N(2 ** i)) mux(
						.data_in(lru_in[(2 ** i) - 1+:2 ** i]),
						.sel_in(tmp[WAY_IDX_BITS - 1-:i]),
						.data_out(tmp[(WAY_IDX_BITS - 1) - i])
					);
				end
			end
			// Trace: src/VX_cache_repl.sv:53:9
			assign way_idx = tmp;
		end
		else begin : g_no_enc
			// Trace: src/VX_cache_repl.sv:55:9
			assign way_idx = 1'sb0;
		end
	endgenerate
endmodule
module VX_cache_repl (
	clk,
	reset,
	stall,
	hit_valid,
	hit_line,
	hit_way,
	repl_valid,
	repl_line,
	repl_way
);
	// Trace: src/VX_cache_repl.sv:59:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_cache_repl.sv:60:15
	parameter LINE_SIZE = 64;
	// Trace: src/VX_cache_repl.sv:61:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_repl.sv:62:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_repl.sv:63:15
	parameter REPL_POLICY = 1;
	// Trace: src/VX_cache_repl.sv:65:5
	input wire clk;
	// Trace: src/VX_cache_repl.sv:66:5
	input wire reset;
	// Trace: src/VX_cache_repl.sv:67:5
	input wire stall;
	// Trace: src/VX_cache_repl.sv:68:5
	input wire hit_valid;
	// Trace: src/VX_cache_repl.sv:69:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] hit_line;
	// Trace: src/VX_cache_repl.sv:70:5
	input wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] hit_way;
	// Trace: src/VX_cache_repl.sv:71:5
	input wire repl_valid;
	// Trace: src/VX_cache_repl.sv:72:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] repl_line;
	// Trace: src/VX_cache_repl.sv:73:5
	output wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] repl_way;
	// Trace: src/VX_cache_repl.sv:75:5
	localparam WAY_SEL_WIDTH = ($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1);
	// Trace: src/VX_cache_repl.sv:76:5
	generate
		if (NUM_WAYS > 1) begin : g_enable
			if (REPL_POLICY == 2) begin : g_plru
				// Trace: src/VX_cache_repl.sv:78:13
				localparam LRU_WIDTH = ((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1);
				// Trace: src/VX_cache_repl.sv:79:13
				wire [LRU_WIDTH - 1:0] plru_rdata;
				// Trace: src/VX_cache_repl.sv:80:13
				wire [LRU_WIDTH - 1:0] plru_wdata;
				// Trace: src/VX_cache_repl.sv:81:13
				wire [LRU_WIDTH - 1:0] plru_wmask;
				// Trace: src/VX_cache_repl.sv:82:13
				VX_dp_ram #(
					.DATAW(LRU_WIDTH),
					.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
					.WRENW(LRU_WIDTH),
					.RDW_MODE("R"),
					.RADDR_REG(1)
				) plru_store(
					.clk(clk),
					.reset(reset),
					.read(repl_valid),
					.write(hit_valid),
					.wren(plru_wmask),
					.waddr(hit_line),
					.raddr(repl_line),
					.wdata(plru_wdata),
					.rdata(plru_rdata)
				);
				// Trace: src/VX_cache_repl.sv:99:13
				plru_decoder #(.NUM_WAYS(NUM_WAYS)) plru_dec(
					.way_idx(hit_way),
					.lru_data(plru_wdata),
					.lru_mask(plru_wmask)
				);
				// Trace: src/VX_cache_repl.sv:106:13
				plru_encoder #(.NUM_WAYS(NUM_WAYS)) plru_enc(
					.lru_in(plru_rdata),
					.way_idx(repl_way)
				);
			end
			else if (REPL_POLICY == 1) begin : g_cyclic
				// Trace: src/VX_cache_repl.sv:113:13
				wire [WAY_SEL_WIDTH - 1:0] ctr_rdata;
				// Trace: src/VX_cache_repl.sv:114:13
				wire [WAY_SEL_WIDTH - 1:0] ctr_wdata = ctr_rdata + 1;
				// Trace: src/VX_cache_repl.sv:115:13
				VX_sp_ram #(
					.DATAW(WAY_SEL_WIDTH),
					.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
					.RDW_MODE("R"),
					.RADDR_REG(1)
				) ctr_store(
					.clk(clk),
					.reset(reset),
					.read(repl_valid),
					.write(repl_valid),
					.wren(1'b1),
					.addr(repl_line),
					.wdata(ctr_wdata),
					.rdata(ctr_rdata)
				);
				// Trace: src/VX_cache_repl.sv:130:13
				assign repl_way = ctr_rdata;
			end
			else begin : g_random
				// Trace: src/VX_cache_repl.sv:132:13
				reg [WAY_SEL_WIDTH - 1:0] victim_idx;
				// Trace: src/VX_cache_repl.sv:133:13
				always @(posedge clk)
					// Trace: src/VX_cache_repl.sv:134:17
					if (reset)
						// Trace: src/VX_cache_repl.sv:135:21
						victim_idx <= 0;
					else if (~stall)
						// Trace: src/VX_cache_repl.sv:137:21
						victim_idx <= victim_idx + 1;
				// Trace: src/VX_cache_repl.sv:140:13
				assign repl_way = victim_idx;
			end
		end
		else begin : g_disable
			// Trace: src/VX_cache_repl.sv:143:9
			assign repl_way = 1'b0;
		end
	endgenerate
endmodule
module VX_stream_omega (
	clk,
	reset,
	valid_in,
	data_in,
	sel_in,
	ready_in,
	valid_out,
	data_out,
	sel_out,
	ready_out,
	collisions
);
	// Trace: src/VX_stream_omega.sv:2:15
	parameter NUM_INPUTS = 4;
	// Trace: src/VX_stream_omega.sv:3:15
	parameter NUM_OUTPUTS = 4;
	// Trace: src/VX_stream_omega.sv:4:15
	parameter RADIX = 2;
	// Trace: src/VX_stream_omega.sv:5:15
	parameter DATAW = 4;
	// Trace: src/VX_stream_omega.sv:6:15
	parameter ARBITER = "R";
	// Trace: src/VX_stream_omega.sv:7:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_omega.sv:8:15
	parameter MAX_FANOUT = 8;
	// Trace: src/VX_stream_omega.sv:9:15
	parameter PERF_CTR_BITS = 32;
	// Trace: src/VX_stream_omega.sv:10:15
	parameter IN_WIDTH = (NUM_INPUTS > 1 ? $clog2(NUM_INPUTS) : 1);
	// Trace: src/VX_stream_omega.sv:11:15
	parameter OUT_WIDTH = (NUM_OUTPUTS > 1 ? $clog2(NUM_OUTPUTS) : 1);
	// Trace: src/VX_stream_omega.sv:13:5
	input wire clk;
	// Trace: src/VX_stream_omega.sv:14:5
	input wire reset;
	// Trace: src/VX_stream_omega.sv:15:5
	input wire [NUM_INPUTS - 1:0] valid_in;
	// Trace: src/VX_stream_omega.sv:16:5
	input wire [(NUM_INPUTS * DATAW) - 1:0] data_in;
	// Trace: src/VX_stream_omega.sv:17:5
	input wire [(NUM_INPUTS * OUT_WIDTH) - 1:0] sel_in;
	// Trace: src/VX_stream_omega.sv:18:5
	output wire [NUM_INPUTS - 1:0] ready_in;
	// Trace: src/VX_stream_omega.sv:19:5
	output wire [NUM_OUTPUTS - 1:0] valid_out;
	// Trace: src/VX_stream_omega.sv:20:5
	output wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out;
	// Trace: src/VX_stream_omega.sv:21:5
	output wire [(NUM_OUTPUTS * IN_WIDTH) - 1:0] sel_out;
	// Trace: src/VX_stream_omega.sv:22:5
	input wire [NUM_OUTPUTS - 1:0] ready_out;
	// Trace: src/VX_stream_omega.sv:23:5
	output wire [PERF_CTR_BITS - 1:0] collisions;
	// Trace: src/VX_stream_omega.sv:25:5
	function automatic [DATAW - 1:0] sv2v_cast_8E21C;
		input reg [DATAW - 1:0] inp;
		sv2v_cast_8E21C = inp;
	endfunction
	function automatic signed [IN_WIDTH - 1:0] sv2v_cast_314B8_signed;
		input reg signed [IN_WIDTH - 1:0] inp;
		sv2v_cast_314B8_signed = inp;
	endfunction
	function automatic [IN_WIDTH - 1:0] sv2v_cast_314B8;
		input reg [IN_WIDTH - 1:0] inp;
		sv2v_cast_314B8 = inp;
	endfunction
	function automatic [PERF_CTR_BITS - 1:0] sv2v_cast_8BEE5;
		input reg [PERF_CTR_BITS - 1:0] inp;
		sv2v_cast_8BEE5 = inp;
	endfunction
	generate
		if ((NUM_INPUTS <= RADIX) && (NUM_OUTPUTS <= RADIX)) begin : g_fallback
			// Trace: src/VX_stream_omega.sv:26:9
			VX_stream_xbar #(
				.NUM_INPUTS(NUM_INPUTS),
				.NUM_OUTPUTS(NUM_OUTPUTS),
				.DATAW(DATAW),
				.ARBITER(ARBITER),
				.OUT_BUF(OUT_BUF),
				.MAX_FANOUT(MAX_FANOUT),
				.PERF_CTR_BITS(PERF_CTR_BITS)
			) xbar_switch(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_in),
				.data_in(data_in),
				.sel_in(sel_in),
				.ready_in(ready_in),
				.valid_out(valid_out),
				.data_out(data_out),
				.sel_out(sel_out),
				.ready_out(ready_out),
				.collisions(collisions)
			);
		end
		else begin : g_omega
			// Trace: src/VX_stream_omega.sv:48:9
			localparam RADIX_LG = (RADIX > 1 ? $clog2(RADIX) : 1);
			// Trace: src/VX_stream_omega.sv:49:9
			localparam N_INPUTS_M = (NUM_INPUTS > NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
			// Trace: src/VX_stream_omega.sv:50:9
			localparam N_INPUTS_LG = (($clog2(N_INPUTS_M) + RADIX_LG) - 1) / RADIX_LG;
			// Trace: src/VX_stream_omega.sv:51:9
			localparam N_INPUTS = RADIX ** N_INPUTS_LG;
			// Trace: src/VX_stream_omega.sv:52:9
			localparam NUM_STAGES = (N_INPUTS > 1 ? $clog2(N_INPUTS) : 1) / RADIX_LG;
			// Trace: src/VX_stream_omega.sv:53:9
			localparam NUM_SWITCHES = N_INPUTS / RADIX;
			// Trace: src/VX_stream_omega.sv:54:9
			// removed localparam type omega_t
			// Trace: src/VX_stream_omega.sv:59:9
			wire [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] switch_valid_in;
			wire [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] switch_valid_out;
			// Trace: src/VX_stream_omega.sv:60:9
			wire [(((NUM_STAGES * NUM_SWITCHES) * RADIX) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) - 1:0] switch_data_in;
			wire [(((NUM_STAGES * NUM_SWITCHES) * RADIX) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) - 1:0] switch_data_out;
			// Trace: src/VX_stream_omega.sv:61:9
			wire [(((NUM_STAGES * NUM_SWITCHES) * RADIX) * RADIX_LG) - 1:0] switch_sel_in;
			// Trace: src/VX_stream_omega.sv:62:9
			wire [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] switch_ready_in;
			wire [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] switch_ready_out;
			genvar _gv_i_3;
			for (_gv_i_3 = 0; _gv_i_3 < N_INPUTS; _gv_i_3 = _gv_i_3 + 1) begin : g_tie_inputs
				localparam i = _gv_i_3;
				// Trace: src/VX_stream_omega.sv:64:13
				localparam DST_IDX = ((i << 1) | (i >> (N_INPUTS_LG - 1))) & (N_INPUTS - 1);
				// Trace: src/VX_stream_omega.sv:65:13
				localparam switch = DST_IDX / RADIX;
				// Trace: src/VX_stream_omega.sv:66:13
				localparam port = DST_IDX % RADIX;
				if (i < NUM_INPUTS) begin : g_valid
					// Trace: src/VX_stream_omega.sv:68:17
					assign switch_valid_in[((0 + switch) * RADIX) + port] = valid_in[i];
					// Trace: src/VX_stream_omega.sv:69:17
					function automatic [N_INPUTS_LG - 1:0] sv2v_cast_51E45;
						input reg [N_INPUTS_LG - 1:0] inp;
						sv2v_cast_51E45 = inp;
					endfunction
					function automatic [N_INPUTS_LG - 1:0] sv2v_cast_43513;
						input reg [N_INPUTS_LG - 1:0] inp;
						sv2v_cast_43513 = inp;
					endfunction
					assign switch_data_in[(((0 + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)+:(N_INPUTS_LG + DATAW) + IN_WIDTH] = {sv2v_cast_43513(sv2v_cast_51E45(sel_in[i * OUT_WIDTH+:OUT_WIDTH])), sv2v_cast_8E21C(data_in[i * DATAW+:DATAW]), sv2v_cast_314B8(sv2v_cast_314B8_signed(i))};
					// Trace: src/VX_stream_omega.sv:74:17
					assign ready_in[i] = switch_ready_in[((0 + switch) * RADIX) + port];
				end
				else begin : g_padding
					// Trace: src/VX_stream_omega.sv:76:17
					assign switch_valid_in[((0 + switch) * RADIX) + port] = 0;
					// Trace: src/VX_stream_omega.sv:77:17
					assign switch_data_in[(((0 + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)+:(N_INPUTS_LG + DATAW) + IN_WIDTH] = 1'sbx;
				end
			end
			genvar _gv_stage_1;
			for (_gv_stage_1 = 0; _gv_stage_1 < NUM_STAGES; _gv_stage_1 = _gv_stage_1 + 1) begin : g_sel_in
				localparam stage = _gv_stage_1;
				genvar _gv_switch_1;
				for (_gv_switch_1 = 0; _gv_switch_1 < NUM_SWITCHES; _gv_switch_1 = _gv_switch_1 + 1) begin : g_switches
					localparam switch = _gv_switch_1;
					genvar _gv_port_1;
					for (_gv_port_1 = 0; _gv_port_1 < RADIX; _gv_port_1 = _gv_port_1 + 1) begin : g_ports
						localparam port = _gv_port_1;
						// Trace: src/VX_stream_omega.sv:83:21
						assign switch_sel_in[((((stage * NUM_SWITCHES) + switch) * RADIX) + port) * RADIX_LG+:RADIX_LG] = switch_data_in[(((((stage * NUM_SWITCHES) + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) + ((N_INPUTS_LG + (DATAW + (IN_WIDTH - 1))) - ((N_INPUTS_LG - 1) - (((NUM_STAGES - 1) - stage) * RADIX_LG)))+:RADIX_LG];
					end
				end
			end
			genvar _gv_stage_2;
			for (_gv_stage_2 = 0; _gv_stage_2 < (NUM_STAGES - 1); _gv_stage_2 = _gv_stage_2 + 1) begin : g_stages
				localparam stage = _gv_stage_2;
				genvar _gv_switch_2;
				for (_gv_switch_2 = 0; _gv_switch_2 < NUM_SWITCHES; _gv_switch_2 = _gv_switch_2 + 1) begin : g_switches
					localparam switch = _gv_switch_2;
					genvar _gv_port_2;
					for (_gv_port_2 = 0; _gv_port_2 < RADIX; _gv_port_2 = _gv_port_2 + 1) begin : g_ports
						localparam port = _gv_port_2;
						// Trace: src/VX_stream_omega.sv:90:21
						localparam lane = (switch * RADIX) + port;
						// Trace: src/VX_stream_omega.sv:91:21
						localparam dst_lane = ((lane << 1) | (lane >> (N_INPUTS_LG - 1))) & (N_INPUTS - 1);
						// Trace: src/VX_stream_omega.sv:92:21
						localparam dst_switch = dst_lane / RADIX;
						// Trace: src/VX_stream_omega.sv:93:21
						localparam dst_port = dst_lane % RADIX;
						// Trace: src/VX_stream_omega.sv:94:21
						assign switch_valid_in[((((stage + 1) * NUM_SWITCHES) + dst_switch) * RADIX) + dst_port] = switch_valid_out[(((stage * NUM_SWITCHES) + switch) * RADIX) + port];
						// Trace: src/VX_stream_omega.sv:95:21
						assign switch_data_in[(((((stage + 1) * NUM_SWITCHES) + dst_switch) * RADIX) + dst_port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)+:(N_INPUTS_LG + DATAW) + IN_WIDTH] = switch_data_out[((((stage * NUM_SWITCHES) + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)+:(N_INPUTS_LG + DATAW) + IN_WIDTH];
						// Trace: src/VX_stream_omega.sv:96:21
						assign switch_ready_out[(((stage * NUM_SWITCHES) + switch) * RADIX) + port] = switch_ready_in[((((stage + 1) * NUM_SWITCHES) + dst_switch) * RADIX) + dst_port];
					end
				end
			end
			genvar _gv_switch_3;
			for (_gv_switch_3 = 0; _gv_switch_3 < NUM_SWITCHES; _gv_switch_3 = _gv_switch_3 + 1) begin : g_switches
				localparam switch = _gv_switch_3;
				genvar _gv_stage_3;
				for (_gv_stage_3 = 0; _gv_stage_3 < NUM_STAGES; _gv_stage_3 = _gv_stage_3 + 1) begin : g_stages
					localparam stage = _gv_stage_3;
					// Trace: src/VX_stream_omega.sv:102:17
					VX_stream_xbar #(
						.NUM_INPUTS(RADIX),
						.NUM_OUTPUTS(RADIX),
						.DATAW((N_INPUTS_LG + DATAW) + IN_WIDTH),
						.ARBITER(ARBITER),
						.OUT_BUF(OUT_BUF),
						.MAX_FANOUT(MAX_FANOUT),
						.PERF_CTR_BITS(PERF_CTR_BITS)
					) xbar_switch(
						.clk(clk),
						.reset(reset),
						.valid_in(switch_valid_in[((stage * NUM_SWITCHES) + switch) * RADIX+:RADIX]),
						.data_in(switch_data_in[((N_INPUTS_LG + DATAW) + IN_WIDTH) * (((stage * NUM_SWITCHES) + switch) * RADIX)+:((N_INPUTS_LG + DATAW) + IN_WIDTH) * RADIX]),
						.sel_in(switch_sel_in[RADIX_LG * (((stage * NUM_SWITCHES) + switch) * RADIX)+:RADIX_LG * RADIX]),
						.ready_in(switch_ready_in[((stage * NUM_SWITCHES) + switch) * RADIX+:RADIX]),
						.valid_out(switch_valid_out[((stage * NUM_SWITCHES) + switch) * RADIX+:RADIX]),
						.data_out(switch_data_out[((N_INPUTS_LG + DATAW) + IN_WIDTH) * (((stage * NUM_SWITCHES) + switch) * RADIX)+:((N_INPUTS_LG + DATAW) + IN_WIDTH) * RADIX]),
						.sel_out(),
						.ready_out(switch_ready_out[((stage * NUM_SWITCHES) + switch) * RADIX+:RADIX]),
						.collisions()
					);
				end
			end
			genvar _gv_i_4;
			for (_gv_i_4 = 0; _gv_i_4 < N_INPUTS; _gv_i_4 = _gv_i_4 + 1) begin : g_tie_outputs
				localparam i = _gv_i_4;
				// Trace: src/VX_stream_omega.sv:126:13
				localparam switch = i / RADIX;
				// Trace: src/VX_stream_omega.sv:127:13
				localparam port = i % RADIX;
				if (i < NUM_OUTPUTS) begin : g_valid
					// Trace: src/VX_stream_omega.sv:129:17
					assign valid_out[i] = switch_valid_out[((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port];
					// Trace: src/VX_stream_omega.sv:130:17
					assign data_out[i * DATAW+:DATAW] = switch_data_out[((((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) + (DATAW + (IN_WIDTH - 1))-:((DATAW + (IN_WIDTH - 1)) >= (IN_WIDTH + 0) ? ((DATAW + (IN_WIDTH - 1)) - (IN_WIDTH + 0)) + 1 : ((IN_WIDTH + 0) - (DATAW + (IN_WIDTH - 1))) + 1)];
					// Trace: src/VX_stream_omega.sv:131:17
					assign sel_out[i * IN_WIDTH+:IN_WIDTH] = switch_data_out[((((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) + (IN_WIDTH - 1)-:IN_WIDTH];
					// Trace: src/VX_stream_omega.sv:132:17
					assign switch_ready_out[((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port] = ready_out[i];
				end
				else begin : g_padding
					// Trace: src/VX_stream_omega.sv:134:17
					assign switch_ready_out[((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port] = 0;
				end
			end
			// Trace: src/VX_stream_omega.sv:137:9
			reg [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] per_cycle_collision;
			reg [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] per_cycle_collision_r;
			// Trace: src/VX_stream_omega.sv:138:9
			wire [$clog2(((NUM_STAGES * NUM_SWITCHES) * RADIX) + 1) - 1:0] collision_count;
			// Trace: src/VX_stream_omega.sv:139:9
			reg [PERF_CTR_BITS - 1:0] collisions_r;
			// Trace: src/VX_stream_omega.sv:140:9
			always @(*) begin
				// Trace: src/VX_stream_omega.sv:141:13
				per_cycle_collision = 0;
				// Trace: src/VX_stream_omega.sv:142:13
				begin : sv2v_autoblock_1
					// Trace: src/VX_stream_omega.sv:142:18
					integer stage;
					// Trace: src/VX_stream_omega.sv:142:18
					for (stage = 0; stage < NUM_STAGES; stage = stage + 1)
						begin
							// Trace: src/VX_stream_omega.sv:143:17
							begin : sv2v_autoblock_2
								// Trace: src/VX_stream_omega.sv:143:22
								integer switch;
								// Trace: src/VX_stream_omega.sv:143:22
								for (switch = 0; switch < NUM_SWITCHES; switch = switch + 1)
									begin
										// Trace: src/VX_stream_omega.sv:144:21
										begin : sv2v_autoblock_3
											// Trace: src/VX_stream_omega.sv:144:26
											integer port_a;
											// Trace: src/VX_stream_omega.sv:144:26
											for (port_a = 0; port_a < RADIX; port_a = port_a + 1)
												begin
													// Trace: src/VX_stream_omega.sv:145:25
													begin : sv2v_autoblock_4
														// Trace: src/VX_stream_omega.sv:145:30
														integer port_b;
														// Trace: src/VX_stream_omega.sv:145:30
														for (port_b = port_a + 1; port_b < RADIX; port_b = port_b + 1)
															begin
																// Trace: src/VX_stream_omega.sv:146:29
																per_cycle_collision[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_a] = per_cycle_collision[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_a] | (((switch_valid_in[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_a] && switch_valid_in[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_b]) && (switch_sel_in[((((stage * NUM_SWITCHES) + switch) * RADIX) + port_a) * RADIX_LG+:RADIX_LG] == switch_sel_in[((((stage * NUM_SWITCHES) + switch) * RADIX) + port_b) * RADIX_LG+:RADIX_LG])) && (switch_ready_in[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_a] | switch_ready_in[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_b]));
															end
													end
												end
										end
									end
							end
						end
				end
			end
			// Trace: src/VX_stream_omega.sv:155:5
			// rewrote reg-to-output bindings
			wire [(NUM_STAGES * NUM_SWITCHES) * RADIX:1] sv2v_tmp___per_cycle_collision_r___data_out;
			always @(*) per_cycle_collision_r = sv2v_tmp___per_cycle_collision_r___data_out;
			VX_pipe_register #(
				.DATAW((NUM_STAGES * NUM_SWITCHES) * RADIX),
				.RESETW(0),
				.DEPTH(1)
			) __per_cycle_collision_r__(
				.clk(clk),
				.reset(reset),
				.enable(1'b1),
				.data_in(per_cycle_collision),
				.data_out(sv2v_tmp___per_cycle_collision_r___data_out)
			);
			// Trace: src/VX_stream_omega.sv:166:5
			VX_popcount #(
				.N((NUM_STAGES * NUM_SWITCHES) * RADIX),
				.MODEL(1)
			) __collision_count__(
				.data_in(per_cycle_collision_r),
				.data_out(collision_count)
			);
			// Trace: src/VX_stream_omega.sv:173:9
			always @(posedge clk)
				// Trace: src/VX_stream_omega.sv:174:13
				if (reset)
					// Trace: src/VX_stream_omega.sv:175:17
					collisions_r <= 1'sb0;
				else
					// Trace: src/VX_stream_omega.sv:177:17
					collisions_r <= collisions_r + sv2v_cast_8BEE5(collision_count);
			// Trace: src/VX_stream_omega.sv:180:9
			assign collisions = collisions_r;
		end
	endgenerate
endmodule
// removed interface: VX_commit_csr_if
// removed module with interface ports: VX_fetch
module VX_pipe_buffer (
	clk,
	reset,
	valid_in,
	ready_in,
	data_in,
	data_out,
	ready_out,
	valid_out
);
	// Trace: src/VX_pipe_buffer.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_pipe_buffer.sv:3:15
	parameter RESETW = 0;
	// Trace: src/VX_pipe_buffer.sv:4:15
	parameter DEPTH = 1;
	// Trace: src/VX_pipe_buffer.sv:6:5
	input wire clk;
	// Trace: src/VX_pipe_buffer.sv:7:5
	input wire reset;
	// Trace: src/VX_pipe_buffer.sv:8:5
	input wire valid_in;
	// Trace: src/VX_pipe_buffer.sv:9:5
	output wire ready_in;
	// Trace: src/VX_pipe_buffer.sv:10:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_pipe_buffer.sv:11:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_pipe_buffer.sv:12:5
	input wire ready_out;
	// Trace: src/VX_pipe_buffer.sv:13:5
	output wire valid_out;
	// Trace: src/VX_pipe_buffer.sv:15:5
	generate
		if (DEPTH == 0) begin : g_passthru
			// Trace: src/VX_pipe_buffer.sv:16:9
			assign ready_in = ready_out;
			// Trace: src/VX_pipe_buffer.sv:17:9
			assign valid_out = valid_in;
			// Trace: src/VX_pipe_buffer.sv:18:9
			assign data_out = data_in;
		end
		else begin : g_register
			// Trace: src/VX_pipe_buffer.sv:20:9
			wire [DEPTH:0] valid;
			// Trace: src/VX_pipe_buffer.sv:21:9
			wire ready [0:DEPTH + 0];
			// Trace: src/VX_pipe_buffer.sv:22:9
			wire [(DEPTH >= 0 ? ((DEPTH + 1) * DATAW) - 1 : ((1 - DEPTH) * DATAW) + ((DEPTH * DATAW) - 1)):(DEPTH >= 0 ? 0 : DEPTH * DATAW)] data;
			// Trace: src/VX_pipe_buffer.sv:23:9
			assign valid[0] = valid_in;
			// Trace: src/VX_pipe_buffer.sv:24:9
			assign data[(DEPTH >= 0 ? 0 : DEPTH) * DATAW+:DATAW] = data_in;
			// Trace: src/VX_pipe_buffer.sv:25:9
			assign ready_in = ready[0];
			genvar _gv_i_7;
			for (_gv_i_7 = 0; _gv_i_7 < DEPTH; _gv_i_7 = _gv_i_7 + 1) begin : g_pipe_regs
				localparam i = _gv_i_7;
				// Trace: src/VX_pipe_buffer.sv:27:13
				assign ready[i] = ready[i + 1] || ~valid[i + 1];
				// Trace: src/VX_pipe_buffer.sv:28:13
				VX_pipe_register #(
					.DATAW(1 + DATAW),
					.RESETW(1 + RESETW)
				) pipe_register(
					.clk(clk),
					.reset(reset),
					.enable(ready[i]),
					.data_in({valid[i], data[(DEPTH >= 0 ? i : DEPTH - i) * DATAW+:DATAW]}),
					.data_out({valid[i + 1], data[(DEPTH >= 0 ? i + 1 : DEPTH - (i + 1)) * DATAW+:DATAW]})
				);
			end
			// Trace: src/VX_pipe_buffer.sv:39:9
			assign valid_out = valid[DEPTH];
			// Trace: src/VX_pipe_buffer.sv:40:9
			assign data_out = data[(DEPTH >= 0 ? DEPTH : DEPTH - DEPTH) * DATAW+:DATAW];
			// Trace: src/VX_pipe_buffer.sv:41:9
			assign ready[DEPTH] = ready_out;
		end
	endgenerate
endmodule
// removed package "VX_gpu_pkg"
// removed interface: VX_dcr_bus_if
// removed module with interface ports: VX_issue_slice
// removed module with interface ports: VX_alu_int
// removed module with interface ports: VX_pe_switch
// removed module with interface ports: VX_wctl_unit
// removed interface: VX_decode_if
// removed interface: VX_execute_if
// removed interface: VX_scoreboard_if
// removed module with interface ports: VX_gbar_unit
// removed module with interface ports: VX_cache
// removed module with interface ports: VX_csr_data
module VX_fifo_queue (
	clk,
	reset,
	push,
	pop,
	data_in,
	data_out,
	empty,
	alm_empty,
	full,
	alm_full,
	size
);
	// Trace: src/VX_fifo_queue.sv:2:15
	parameter DATAW = 32;
	// Trace: src/VX_fifo_queue.sv:3:15
	parameter DEPTH = 32;
	// Trace: src/VX_fifo_queue.sv:4:15
	parameter ALM_FULL = DEPTH - 1;
	// Trace: src/VX_fifo_queue.sv:5:15
	parameter ALM_EMPTY = 1;
	// Trace: src/VX_fifo_queue.sv:6:15
	parameter OUT_REG = 0;
	// Trace: src/VX_fifo_queue.sv:7:15
	parameter LUTRAM = 0;
	// Trace: src/VX_fifo_queue.sv:8:15
	parameter SIZEW = $clog2(DEPTH + 1);
	// Trace: src/VX_fifo_queue.sv:10:5
	input wire clk;
	// Trace: src/VX_fifo_queue.sv:11:5
	input wire reset;
	// Trace: src/VX_fifo_queue.sv:12:5
	input wire push;
	// Trace: src/VX_fifo_queue.sv:13:5
	input wire pop;
	// Trace: src/VX_fifo_queue.sv:14:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_fifo_queue.sv:15:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_fifo_queue.sv:16:5
	output wire empty;
	// Trace: src/VX_fifo_queue.sv:17:5
	output wire alm_empty;
	// Trace: src/VX_fifo_queue.sv:18:5
	output wire full;
	// Trace: src/VX_fifo_queue.sv:19:5
	output wire alm_full;
	// Trace: src/VX_fifo_queue.sv:20:5
	output wire [SIZEW - 1:0] size;
	// Trace: src/VX_fifo_queue.sv:22:5
	VX_pending_size #(
		.SIZE(DEPTH),
		.ALM_EMPTY(ALM_EMPTY),
		.ALM_FULL(ALM_FULL)
	) pending_size(
		.clk(clk),
		.reset(reset),
		.incr(push),
		.decr(pop),
		.empty(empty),
		.full(full),
		.alm_empty(alm_empty),
		.alm_full(alm_full),
		.size(size)
	);
	// Trace: src/VX_fifo_queue.sv:37:5
	generate
		if (DEPTH == 1) begin : g_depth_1
			// Trace: src/VX_fifo_queue.sv:38:9
			reg [DATAW - 1:0] head_r;
			// Trace: src/VX_fifo_queue.sv:39:9
			always @(posedge clk)
				// Trace: src/VX_fifo_queue.sv:40:13
				if (push)
					// Trace: src/VX_fifo_queue.sv:41:17
					head_r <= data_in;
			// Trace: src/VX_fifo_queue.sv:44:9
			assign data_out = head_r;
		end
		else begin : g_depth_n
			// Trace: src/VX_fifo_queue.sv:46:9
			localparam ADDRW = $clog2(DEPTH);
			// Trace: src/VX_fifo_queue.sv:47:9
			wire [DATAW - 1:0] data_out_w;
			// Trace: src/VX_fifo_queue.sv:48:9
			reg [ADDRW - 1:0] rd_ptr_r;
			// Trace: src/VX_fifo_queue.sv:49:9
			reg [ADDRW - 1:0] wr_ptr_r;
			// Trace: src/VX_fifo_queue.sv:50:9
			always @(posedge clk)
				// Trace: src/VX_fifo_queue.sv:51:13
				if (reset) begin
					// Trace: src/VX_fifo_queue.sv:52:17
					wr_ptr_r <= 1'sb0;
					// Trace: src/VX_fifo_queue.sv:53:17
					rd_ptr_r <= (OUT_REG != 0 ? 1 : 0);
				end
				else begin
					// Trace: src/VX_fifo_queue.sv:55:17
					begin : sv2v_autoblock_1
						reg [ADDRW - 1:0] sv2v_tmp_cast;
						sv2v_tmp_cast = push;
						wr_ptr_r <= wr_ptr_r + sv2v_tmp_cast;
					end
					// Trace: src/VX_fifo_queue.sv:56:17
					begin : sv2v_autoblock_2
						reg [ADDRW - 1:0] sv2v_tmp_cast_1;
						sv2v_tmp_cast_1 = pop;
						rd_ptr_r <= rd_ptr_r + sv2v_tmp_cast_1;
					end
				end
			// Trace: src/VX_fifo_queue.sv:59:9
			VX_dp_ram #(
				.DATAW(DATAW),
				.SIZE(DEPTH),
				.LUTRAM(LUTRAM),
				.RDW_MODE("W"),
				.RADDR_REG(1)
			) dp_ram(
				.clk(clk),
				.reset(reset),
				.read(1'b1),
				.write(push),
				.wren(1'b1),
				.raddr(rd_ptr_r),
				.waddr(wr_ptr_r),
				.wdata(data_in),
				.rdata(data_out_w)
			);
			if (OUT_REG != 0) begin : g_out_reg
				// Trace: src/VX_fifo_queue.sv:77:13
				reg [DATAW - 1:0] data_out_r;
				// Trace: src/VX_fifo_queue.sv:78:13
				function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
					input reg signed [ADDRW - 1:0] inp;
					sv2v_cast_8BB5D_signed = inp;
				endfunction
				wire going_empty = (ALM_EMPTY == 1 ? alm_empty : size[ADDRW - 1:0] == sv2v_cast_8BB5D_signed(1));
				// Trace: src/VX_fifo_queue.sv:79:13
				wire bypass = push && (empty || (going_empty && pop));
				// Trace: src/VX_fifo_queue.sv:80:13
				always @(posedge clk)
					// Trace: src/VX_fifo_queue.sv:81:17
					if (bypass)
						// Trace: src/VX_fifo_queue.sv:82:21
						data_out_r <= data_in;
					else if (pop)
						// Trace: src/VX_fifo_queue.sv:84:21
						data_out_r <= data_out_w;
				// Trace: src/VX_fifo_queue.sv:87:13
				assign data_out = data_out_r;
			end
			else begin : g_no_out_reg
				// Trace: src/VX_fifo_queue.sv:89:13
				assign data_out = data_out_w;
			end
		end
	endgenerate
endmodule
// removed module with interface ports: VX_commit
module VX_stream_unpack (
	clk,
	reset,
	valid_in,
	mask_in,
	data_in,
	tag_in,
	ready_in,
	valid_out,
	data_out,
	tag_out,
	ready_out
);
	// Trace: src/VX_stream_unpack.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_stream_unpack.sv:3:15
	parameter DATA_WIDTH = 1;
	// Trace: src/VX_stream_unpack.sv:4:15
	parameter TAG_WIDTH = 1;
	// Trace: src/VX_stream_unpack.sv:5:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_unpack.sv:7:5
	input wire clk;
	// Trace: src/VX_stream_unpack.sv:8:5
	input wire reset;
	// Trace: src/VX_stream_unpack.sv:9:5
	input wire valid_in;
	// Trace: src/VX_stream_unpack.sv:10:5
	input wire [NUM_REQS - 1:0] mask_in;
	// Trace: src/VX_stream_unpack.sv:11:5
	input wire [(NUM_REQS * DATA_WIDTH) - 1:0] data_in;
	// Trace: src/VX_stream_unpack.sv:12:5
	input wire [TAG_WIDTH - 1:0] tag_in;
	// Trace: src/VX_stream_unpack.sv:13:5
	output wire ready_in;
	// Trace: src/VX_stream_unpack.sv:14:5
	output wire [NUM_REQS - 1:0] valid_out;
	// Trace: src/VX_stream_unpack.sv:15:5
	output wire [(NUM_REQS * DATA_WIDTH) - 1:0] data_out;
	// Trace: src/VX_stream_unpack.sv:16:5
	output wire [(NUM_REQS * TAG_WIDTH) - 1:0] tag_out;
	// Trace: src/VX_stream_unpack.sv:17:5
	input wire [NUM_REQS - 1:0] ready_out;
	// Trace: src/VX_stream_unpack.sv:19:5
	generate
		if (NUM_REQS > 1) begin : g_unpack
			// Trace: src/VX_stream_unpack.sv:20:9
			reg [NUM_REQS - 1:0] rem_mask_r;
			// Trace: src/VX_stream_unpack.sv:21:9
			wire [NUM_REQS - 1:0] ready_out_w;
			// Trace: src/VX_stream_unpack.sv:22:9
			wire [NUM_REQS - 1:0] rem_mask_n = rem_mask_r & ~ready_out_w;
			// Trace: src/VX_stream_unpack.sv:23:9
			wire sent_all = ~(|(mask_in & rem_mask_n));
			// Trace: src/VX_stream_unpack.sv:24:9
			always @(posedge clk)
				// Trace: src/VX_stream_unpack.sv:25:13
				if (reset)
					// Trace: src/VX_stream_unpack.sv:26:17
					rem_mask_r <= 1'sb1;
				else
					// Trace: src/VX_stream_unpack.sv:28:17
					if (valid_in)
						// Trace: src/VX_stream_unpack.sv:29:21
						rem_mask_r <= (sent_all ? {NUM_REQS {1'sb1}} : rem_mask_n);
			// Trace: src/VX_stream_unpack.sv:33:9
			assign ready_in = sent_all;
			genvar _gv_i_49;
			for (_gv_i_49 = 0; _gv_i_49 < NUM_REQS; _gv_i_49 = _gv_i_49 + 1) begin : g_outbuf
				localparam i = _gv_i_49;
				// Trace: src/VX_stream_unpack.sv:35:13
				VX_elastic_buffer #(
					.DATAW(DATA_WIDTH + TAG_WIDTH),
					.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
					.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
				) out_buf(
					.clk(clk),
					.reset(reset),
					.valid_in((valid_in && mask_in[i]) && rem_mask_r[i]),
					.ready_in(ready_out_w[i]),
					.data_in({data_in[i * DATA_WIDTH+:DATA_WIDTH], tag_in}),
					.data_out({data_out[i * DATA_WIDTH+:DATA_WIDTH], tag_out[i * TAG_WIDTH+:TAG_WIDTH]}),
					.valid_out(valid_out[i]),
					.ready_out(ready_out[i])
				);
			end
		end
		else begin : g_passthru
			// Trace: src/VX_stream_unpack.sv:51:9
			assign valid_out = valid_in;
			// Trace: src/VX_stream_unpack.sv:52:9
			assign data_out = data_in;
			// Trace: src/VX_stream_unpack.sv:53:9
			assign tag_out = tag_in;
			// Trace: src/VX_stream_unpack.sv:54:9
			assign ready_in = ready_out;
		end
	endgenerate
endmodule
// removed interface: VX_decode_sched_if
module VX_fpu_fpnew (
	clk,
	reset,
	valid_in,
	ready_in,
	mask_in,
	tag_in,
	op_type,
	fmt,
	frm,
	dataa,
	datab,
	datac,
	result,
	has_fflags,
	fflags,
	tag_out,
	ready_out,
	valid_out
);
	// removed import VX_fpu_pkg::*;
	// removed import fpnew_pkg::*;
	// removed import cf_math_pkg::*;
	// removed import defs_div_sqrt_mvp::*;
	// Trace: src/VX_fpu_fpnew.sv:7:15
	parameter NUM_LANES = 1;
	// Trace: src/VX_fpu_fpnew.sv:8:15
	parameter TAG_WIDTH = 1;
	// Trace: src/VX_fpu_fpnew.sv:9:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_fpu_fpnew.sv:11:5
	input wire clk;
	// Trace: src/VX_fpu_fpnew.sv:12:5
	input wire reset;
	// Trace: src/VX_fpu_fpnew.sv:13:5
	input wire valid_in;
	// Trace: src/VX_fpu_fpnew.sv:14:5
	output wire ready_in;
	// Trace: src/VX_fpu_fpnew.sv:15:5
	input wire [NUM_LANES - 1:0] mask_in;
	// Trace: src/VX_fpu_fpnew.sv:16:5
	input wire [TAG_WIDTH - 1:0] tag_in;
	// Trace: src/VX_fpu_fpnew.sv:17:5
	input wire [3:0] op_type;
	// Trace: src/VX_fpu_fpnew.sv:18:5
	input wire [1:0] fmt;
	// Trace: src/VX_fpu_fpnew.sv:19:5
	input wire [2:0] frm;
	// Trace: src/VX_fpu_fpnew.sv:20:5
	input wire [(NUM_LANES * 32) - 1:0] dataa;
	// Trace: src/VX_fpu_fpnew.sv:21:5
	input wire [(NUM_LANES * 32) - 1:0] datab;
	// Trace: src/VX_fpu_fpnew.sv:22:5
	input wire [(NUM_LANES * 32) - 1:0] datac;
	// Trace: src/VX_fpu_fpnew.sv:23:5
	output wire [(NUM_LANES * 32) - 1:0] result;
	// Trace: src/VX_fpu_fpnew.sv:24:5
	output wire has_fflags;
	// Trace: src/VX_fpu_fpnew.sv:25:5
	// removed localparam type VX_fpu_pkg_fflags_t
	output wire [4:0] fflags;
	// Trace: src/VX_fpu_fpnew.sv:26:5
	output wire [TAG_WIDTH - 1:0] tag_out;
	// Trace: src/VX_fpu_fpnew.sv:27:5
	input wire ready_out;
	// Trace: src/VX_fpu_fpnew.sv:28:5
	output wire valid_out;
	// Trace: src/VX_fpu_fpnew.sv:30:5
	localparam LATENCY_FDIVSQRT = 16;
	// Trace: src/VX_fpu_fpnew.sv:31:5
	localparam RSP_DATAW = ((NUM_LANES * 32) + 6) + TAG_WIDTH;
	// Trace: src/VX_fpu_fpnew.sv:32:5
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	// removed localparam type fpnew_pkg_fpu_features_t
	localparam [42:0] FPU_FEATURES = {$unsigned(32), 11'b00100000010};
	// Trace: src/VX_fpu_fpnew.sv:39:5
	// removed localparam type fpnew_pkg_pipe_config_t
	// removed localparam type fpnew_pkg_unit_type_t
	localparam [31:0] fpnew_pkg_NUM_OPGROUPS = 4;
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unit_types_t
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unsigned_t
	// removed localparam type fpnew_pkg_fpu_implementation_t
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 32) - 1:0] sv2v_cast_CDC93;
		input reg [((32'd4 * 32'd5) * 32) - 1:0] inp;
		sv2v_cast_CDC93 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 2) - 1:0] sv2v_cast_15FEF;
		input reg [((32'd4 * 32'd5) * 2) - 1:0] inp;
		sv2v_cast_15FEF = inp;
	endfunction
	localparam [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] FPU_IMPLEMENTATION = {sv2v_cast_CDC93({160'h0000000400000000000000000000000000000000, {fpnew_pkg_NUM_FP_FORMATS {sv2v_cast_32($unsigned(LATENCY_FDIVSQRT))}}, {fpnew_pkg_NUM_FP_FORMATS {32'd2}}, {fpnew_pkg_NUM_FP_FORMATS {32'd5}}}), sv2v_cast_15FEF({{fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}, {fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}}), 2'd3};
	// Trace: src/VX_fpu_fpnew.sv:50:5
	wire fpu_ready_in;
	wire fpu_valid_in;
	// Trace: src/VX_fpu_fpnew.sv:51:5
	wire fpu_ready_out;
	wire fpu_valid_out;
	// Trace: src/VX_fpu_fpnew.sv:52:5
	reg [TAG_WIDTH - 1:0] fpu_tag_in;
	reg [TAG_WIDTH - 1:0] fpu_tag_out;
	// Trace: src/VX_fpu_fpnew.sv:53:5
	reg [((3 * NUM_LANES) * 32) - 1:0] fpu_operands;
	// Trace: src/VX_fpu_fpnew.sv:54:5
	wire [(NUM_LANES * 32) - 1:0] fpu_result;
	// Trace: src/VX_fpu_fpnew.sv:55:5
	// removed localparam type fpnew_pkg_status_t
	wire [4:0] fpu_status;
	// Trace: src/VX_fpu_fpnew.sv:56:5
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	reg [3:0] fpu_op;
	// Trace: src/VX_fpu_fpnew.sv:57:5
	reg [2:0] fpu_rnd;
	// Trace: src/VX_fpu_fpnew.sv:58:5
	reg fpu_op_mod;
	// Trace: src/VX_fpu_fpnew.sv:59:5
	reg fpu_has_fflags;
	reg fpu_has_fflags_out;
	// Trace: src/VX_fpu_fpnew.sv:60:5
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	reg [2:0] fpu_src_fmt;
	reg [2:0] fpu_dst_fmt;
	// Trace: src/VX_fpu_fpnew.sv:61:5
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	reg [1:0] fpu_int_fmt;
	// Trace: src/VX_fpu_fpnew.sv:62:5
	function automatic [3:0] sv2v_cast_F1C4D;
		input reg [3:0] inp;
		sv2v_cast_F1C4D = inp;
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	always @(*) begin
		// Trace: src/VX_fpu_fpnew.sv:63:9
		fpu_op = sv2v_cast_F1C4D(1'sbx);
		// Trace: src/VX_fpu_fpnew.sv:64:9
		fpu_rnd = frm;
		// Trace: src/VX_fpu_fpnew.sv:65:9
		fpu_op_mod = 0;
		// Trace: src/VX_fpu_fpnew.sv:66:9
		fpu_has_fflags = 1;
		// Trace: src/VX_fpu_fpnew.sv:67:9
		fpu_operands[0+:32 * NUM_LANES] = dataa;
		// Trace: src/VX_fpu_fpnew.sv:68:9
		fpu_operands[32 * NUM_LANES+:32 * NUM_LANES] = datab;
		// Trace: src/VX_fpu_fpnew.sv:69:9
		fpu_operands[32 * (2 * NUM_LANES)+:32 * NUM_LANES] = datac;
		// Trace: src/VX_fpu_fpnew.sv:70:9
		fpu_dst_fmt = sv2v_cast_0BC43('d0);
		// Trace: src/VX_fpu_fpnew.sv:71:9
		fpu_int_fmt = sv2v_cast_87CC5(2);
		// Trace: src/VX_fpu_fpnew.sv:72:9
		fpu_src_fmt = fpu_dst_fmt;
		// Trace: src/VX_fpu_fpnew.sv:73:9
		case (op_type)
			4'b0000: begin
				// Trace: src/VX_fpu_fpnew.sv:75:17
				fpu_op = sv2v_cast_A53F3(2);
				// Trace: src/VX_fpu_fpnew.sv:76:17
				fpu_operands[32 * NUM_LANES+:32 * NUM_LANES] = dataa;
				// Trace: src/VX_fpu_fpnew.sv:77:17
				fpu_operands[32 * (2 * NUM_LANES)+:32 * NUM_LANES] = datab;
				// Trace: src/VX_fpu_fpnew.sv:78:17
				fpu_op_mod = fmt[1];
			end
			4'b0001:
				// Trace: src/VX_fpu_fpnew.sv:80:30
				fpu_op = sv2v_cast_A53F3(3);
			4'b0010: begin
				// Trace: src/VX_fpu_fpnew.sv:81:29
				fpu_op = sv2v_cast_A53F3(0);
				// Trace: src/VX_fpu_fpnew.sv:81:56
				fpu_op_mod = fmt[1];
			end
			4'b0011: begin
				// Trace: src/VX_fpu_fpnew.sv:82:28
				fpu_op = sv2v_cast_A53F3(1);
				// Trace: src/VX_fpu_fpnew.sv:82:56
				fpu_op_mod = ~fmt[1];
			end
			4'b0100:
				// Trace: src/VX_fpu_fpnew.sv:83:30
				fpu_op = sv2v_cast_A53F3(4);
			4'b0101:
				// Trace: src/VX_fpu_fpnew.sv:84:29
				fpu_op = sv2v_cast_A53F3(5);
			4'b1000, 4'b1001: begin
				// Trace: src/VX_fpu_fpnew.sv:86:28
				fpu_op = sv2v_cast_A53F3(11);
				// Trace: src/VX_fpu_fpnew.sv:86:53
				fpu_op_mod = op_type[0];
			end
			4'b1010, 4'b1011: begin
				// Trace: src/VX_fpu_fpnew.sv:88:28
				fpu_op = sv2v_cast_A53F3(12);
				// Trace: src/VX_fpu_fpnew.sv:88:53
				fpu_op_mod = op_type[0];
			end
			4'b1100:
				// Trace: src/VX_fpu_fpnew.sv:89:28
				fpu_op = sv2v_cast_A53F3(8);
			4'b1110:
				// Trace: src/VX_fpu_fpnew.sv:91:17
				case (frm)
					0, 1, 2: begin
						// Trace: src/VX_fpu_fpnew.sv:92:34
						fpu_op = sv2v_cast_A53F3(6);
						// Trace: src/VX_fpu_fpnew.sv:92:60
						fpu_rnd = {1'b0, frm[1:0]};
						// Trace: src/VX_fpu_fpnew.sv:92:88
						fpu_has_fflags = 0;
					end
					3: begin
						// Trace: src/VX_fpu_fpnew.sv:93:34
						fpu_op = sv2v_cast_A53F3(9);
						// Trace: src/VX_fpu_fpnew.sv:93:64
						fpu_has_fflags = 0;
					end
					4, 5: begin
						// Trace: src/VX_fpu_fpnew.sv:94:34
						fpu_op = sv2v_cast_A53F3(6);
						// Trace: src/VX_fpu_fpnew.sv:94:60
						fpu_rnd = 3'b011;
						// Trace: src/VX_fpu_fpnew.sv:94:78
						fpu_op_mod = ~frm[0];
						// Trace: src/VX_fpu_fpnew.sv:94:100
						fpu_has_fflags = 0;
					end
					6, 7: begin
						// Trace: src/VX_fpu_fpnew.sv:95:34
						fpu_op = sv2v_cast_A53F3(7);
						// Trace: src/VX_fpu_fpnew.sv:95:62
						fpu_rnd = {2'b00, frm[0]};
					end
				endcase
			default:
				;
		endcase
	end
	// Trace: src/VX_fpu_fpnew.sv:101:5
	genvar _gv_i_50;
	// removed localparam type fpnew_pkg_divsqrt_unit_t
	// removed localparam type fpnew_pkg_roundmode_e
	generate
		for (_gv_i_50 = 0; _gv_i_50 < NUM_LANES; _gv_i_50 = _gv_i_50 + 1) begin : g_fpnew_coreses
			localparam i = _gv_i_50;
			// Trace: src/VX_fpu_fpnew.sv:102:9
			wire [TAG_WIDTH + 0:0] fpu_tag;
			// Trace: src/VX_fpu_fpnew.sv:103:9
			wire fpu_valid_out_uq;
			// Trace: src/VX_fpu_fpnew.sv:104:9
			wire fpu_ready_in_uq;
			// Trace: src/VX_fpu_fpnew.sv:105:9
			wire [4:0] fpu_status_uq;
			// Trace: src/VX_fpu_fpnew.sv:106:9
			fpnew_top_7C2B2_D4A54 #(
				.TagType_TAG_WIDTH(TAG_WIDTH),
				.Features(FPU_FEATURES),
				.Implementation(FPU_IMPLEMENTATION),
				.DivSqrtSel(2'd0)
			) fpnew_core(
				.clk_i(clk),
				.rst_ni(~reset),
				.operands_i({fpu_operands[((2 * NUM_LANES) + i) * 32+:32], fpu_operands[(NUM_LANES + i) * 32+:32], fpu_operands[(0 + i) * 32+:32]}),
				.rnd_mode_i(fpu_rnd),
				.op_i(fpu_op),
				.op_mod_i(fpu_op_mod),
				.src_fmt_i(fpu_src_fmt),
				.dst_fmt_i(fpu_dst_fmt),
				.int_fmt_i(fpu_int_fmt),
				.vectorial_op_i(1'b0),
				.simd_mask_i(1'b1),
				.tag_i({fpu_tag_in, fpu_has_fflags}),
				.in_valid_i(fpu_valid_in),
				.in_ready_o(fpu_ready_in_uq),
				.flush_i(1'b0),
				.result_o(fpu_result[i * 32+:32]),
				.status_o(fpu_status_uq),
				.tag_o(fpu_tag),
				.out_valid_o(fpu_valid_out_uq),
				.out_ready_i(fpu_ready_out),
				.busy_o()
			);
			if (i == 0) begin : g_output_0
				// Trace: src/VX_fpu_fpnew.sv:135:13
				wire [(0 + TAG_WIDTH) + 1:1] sv2v_tmp_65428;
				assign sv2v_tmp_65428 = fpu_tag;
				always @(*) {fpu_tag_out, fpu_has_fflags_out} = sv2v_tmp_65428;
				// Trace: src/VX_fpu_fpnew.sv:136:13
				assign fpu_valid_out = fpu_valid_out_uq;
				// Trace: src/VX_fpu_fpnew.sv:137:13
				assign fpu_ready_in = fpu_ready_in_uq;
				// Trace: src/VX_fpu_fpnew.sv:138:13
				assign fpu_status = fpu_status_uq;
			end
		end
	endgenerate
	// Trace: src/VX_fpu_fpnew.sv:141:5
	assign fpu_valid_in = valid_in;
	// Trace: src/VX_fpu_fpnew.sv:142:5
	assign ready_in = fpu_ready_in;
	// Trace: src/VX_fpu_fpnew.sv:143:5
	wire [TAG_WIDTH:1] sv2v_tmp_14562;
	assign sv2v_tmp_14562 = tag_in;
	always @(*) fpu_tag_in = sv2v_tmp_14562;
	// Trace: src/VX_fpu_fpnew.sv:144:5
	VX_elastic_buffer #(
		.DATAW(RSP_DATAW),
		.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
		.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
	) rsp_buf(
		.clk(clk),
		.reset(reset),
		.valid_in(fpu_valid_out),
		.ready_in(fpu_ready_out),
		.data_in({fpu_result, fpu_has_fflags_out, fpu_status, fpu_tag_out}),
		.data_out({result, has_fflags, fflags, tag_out}),
		.valid_out(valid_out),
		.ready_out(ready_out)
	);
endmodule
// removed interface: VX_sched_csr_if
module VX_stream_buffer (
	clk,
	reset,
	valid_in,
	ready_in,
	data_in,
	data_out,
	ready_out,
	valid_out
);
	// Trace: src/VX_stream_buffer.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_stream_buffer.sv:3:12
	parameter OUT_REG = 0;
	// Trace: src/VX_stream_buffer.sv:4:15
	parameter PASSTHRU = 0;
	// Trace: src/VX_stream_buffer.sv:6:5
	input wire clk;
	// Trace: src/VX_stream_buffer.sv:7:5
	input wire reset;
	// Trace: src/VX_stream_buffer.sv:8:5
	input wire valid_in;
	// Trace: src/VX_stream_buffer.sv:9:5
	output wire ready_in;
	// Trace: src/VX_stream_buffer.sv:10:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_stream_buffer.sv:11:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_stream_buffer.sv:12:5
	input wire ready_out;
	// Trace: src/VX_stream_buffer.sv:13:5
	output wire valid_out;
	// Trace: src/VX_stream_buffer.sv:15:5
	generate
		if (PASSTHRU != 0) begin : g_passthru
			// Trace: src/VX_stream_buffer.sv:16:9
			assign ready_in = ready_out;
			// Trace: src/VX_stream_buffer.sv:17:9
			assign valid_out = valid_in;
			// Trace: src/VX_stream_buffer.sv:18:9
			assign data_out = data_in;
		end
		else begin : g_buffer
			// Trace: src/VX_stream_buffer.sv:20:3
			reg [DATAW - 1:0] data_out_r;
			reg [DATAW - 1:0] buffer_r;
			// Trace: src/VX_stream_buffer.sv:21:3
			reg valid_out_r;
			reg valid_in_r;
			// Trace: src/VX_stream_buffer.sv:22:3
			wire fire_in = valid_in && ready_in;
			// Trace: src/VX_stream_buffer.sv:23:3
			wire flow_out = ready_out || ~valid_out;
			// Trace: src/VX_stream_buffer.sv:24:3
			always @(posedge clk)
				// Trace: src/VX_stream_buffer.sv:25:4
				if (reset)
					// Trace: src/VX_stream_buffer.sv:26:5
					valid_in_r <= 1'b1;
				else if (valid_in || flow_out)
					// Trace: src/VX_stream_buffer.sv:28:5
					valid_in_r <= flow_out;
			// Trace: src/VX_stream_buffer.sv:31:3
			always @(posedge clk)
				// Trace: src/VX_stream_buffer.sv:32:4
				if (reset)
					// Trace: src/VX_stream_buffer.sv:33:5
					valid_out_r <= 1'b0;
				else if (flow_out)
					// Trace: src/VX_stream_buffer.sv:35:5
					valid_out_r <= valid_in || ~valid_in_r;
			if (OUT_REG != 0) begin : g_out_reg
				// Trace: src/VX_stream_buffer.sv:39:4
				always @(posedge clk)
					// Trace: src/VX_stream_buffer.sv:40:5
					if (fire_in)
						// Trace: src/VX_stream_buffer.sv:41:6
						buffer_r <= data_in;
				// Trace: src/VX_stream_buffer.sv:44:4
				always @(posedge clk)
					// Trace: src/VX_stream_buffer.sv:45:5
					if (flow_out)
						// Trace: src/VX_stream_buffer.sv:46:6
						data_out_r <= (valid_in_r ? data_in : buffer_r);
				// Trace: src/VX_stream_buffer.sv:49:4
				assign data_out = data_out_r;
			end
			else begin : g_no_out_reg
				// Trace: src/VX_stream_buffer.sv:51:4
				always @(posedge clk)
					// Trace: src/VX_stream_buffer.sv:52:5
					if (fire_in)
						// Trace: src/VX_stream_buffer.sv:53:6
						data_out_r <= data_in;
				// Trace: src/VX_stream_buffer.sv:56:4
				always @(posedge clk)
					// Trace: src/VX_stream_buffer.sv:57:5
					if (fire_in)
						// Trace: src/VX_stream_buffer.sv:58:6
						buffer_r <= data_out_r;
				// Trace: src/VX_stream_buffer.sv:61:4
				assign data_out = (valid_in_r ? data_out_r : buffer_r);
			end
			// Trace: src/VX_stream_buffer.sv:63:3
			assign valid_out = valid_out_r;
			// Trace: src/VX_stream_buffer.sv:64:3
			assign ready_in = valid_in_r;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_issue
// removed module with interface ports: VX_lsu_slice
module VX_generic_arbiter (
	clk,
	reset,
	requests,
	grant_index,
	grant_onehot,
	grant_valid,
	grant_ready
);
	// Trace: src/VX_generic_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_generic_arbiter.sv:3:15
	parameter TYPE = "P";
	// Trace: src/VX_generic_arbiter.sv:4:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_generic_arbiter.sv:6:5
	input wire clk;
	// Trace: src/VX_generic_arbiter.sv:7:5
	input wire reset;
	// Trace: src/VX_generic_arbiter.sv:8:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_generic_arbiter.sv:9:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_generic_arbiter.sv:10:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_generic_arbiter.sv:11:5
	output wire grant_valid;
	// Trace: src/VX_generic_arbiter.sv:12:5
	input wire grant_ready;
	// Trace: src/VX_generic_arbiter.sv:14:5
	generate
		if (TYPE == "P") begin : g_priority
			// Trace: src/VX_generic_arbiter.sv:15:9
			VX_priority_arbiter #(.NUM_REQS(NUM_REQS)) priority_arbiter(
				.requests(requests),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(grant_onehot)
			);
		end
		else if (TYPE == "R") begin : g_round_robin
			// Trace: src/VX_generic_arbiter.sv:24:9
			VX_rr_arbiter #(.NUM_REQS(NUM_REQS)) rr_arbiter(
				.clk(clk),
				.reset(reset),
				.requests(requests),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(grant_onehot),
				.grant_ready(grant_ready)
			);
		end
		else if (TYPE == "M") begin : g_matrix
			// Trace: src/VX_generic_arbiter.sv:36:9
			VX_matrix_arbiter #(.NUM_REQS(NUM_REQS)) matrix_arbiter(
				.clk(clk),
				.reset(reset),
				.requests(requests),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(grant_onehot),
				.grant_ready(grant_ready)
			);
		end
		else if (TYPE == "C") begin : g_cyclic
			// Trace: src/VX_generic_arbiter.sv:48:9
			VX_cyclic_arbiter #(.NUM_REQS(NUM_REQS)) cyclic_arbiter(
				.clk(clk),
				.reset(reset),
				.requests(requests),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(grant_onehot),
				.grant_ready(grant_ready)
			);
		end
	endgenerate
endmodule
// removed interface: VX_schedule_if
module VX_lzc (
	data_in,
	data_out,
	valid_out
);
	// Trace: src/VX_lzc.sv:2:15
	parameter N = 2;
	// Trace: src/VX_lzc.sv:3:15
	parameter REVERSE = 0;
	// Trace: src/VX_lzc.sv:4:15
	parameter LOGN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_lzc.sv:6:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_lzc.sv:7:5
	output wire [LOGN - 1:0] data_out;
	// Trace: src/VX_lzc.sv:8:5
	output wire valid_out;
	// Trace: src/VX_lzc.sv:10:5
	function automatic signed [LOGN - 1:0] sv2v_cast_B9644_signed;
		input reg signed [LOGN - 1:0] inp;
		sv2v_cast_B9644_signed = inp;
	endfunction
	generate
		if (N == 1) begin : g_passthru
			// Trace: src/VX_lzc.sv:11:9
			assign data_out = 1'sb0;
			// Trace: src/VX_lzc.sv:12:9
			assign valid_out = data_in;
		end
		else begin : g_lzc
			// Trace: src/VX_lzc.sv:14:9
			wire [(N * LOGN) - 1:0] indices;
			genvar _gv_i_64;
			for (_gv_i_64 = 0; _gv_i_64 < N; _gv_i_64 = _gv_i_64 + 1) begin : g_indices
				localparam i = _gv_i_64;
				// Trace: src/VX_lzc.sv:16:13
				assign indices[i * LOGN+:LOGN] = (REVERSE ? sv2v_cast_B9644_signed(i) : sv2v_cast_B9644_signed((N - 1) - i));
			end
			// Trace: src/VX_lzc.sv:18:9
			VX_find_first #(
				.N(N),
				.DATAW(LOGN),
				.REVERSE(!REVERSE)
			) find_first(
				.data_in(indices),
				.valid_in(data_in),
				.data_out(data_out),
				.valid_out(valid_out)
			);
		end
	endgenerate
endmodule
// removed interface: VX_pipeline_perf_if
// removed interface: VX_fetch_if
// removed module with interface ports: VX_cache_cluster
module VX_stream_xbar (
	clk,
	reset,
	valid_in,
	data_in,
	sel_in,
	ready_in,
	valid_out,
	data_out,
	sel_out,
	ready_out,
	collisions
);
	// Trace: src/VX_stream_xbar.sv:2:15
	parameter NUM_INPUTS = 4;
	// Trace: src/VX_stream_xbar.sv:3:15
	parameter NUM_OUTPUTS = 4;
	// Trace: src/VX_stream_xbar.sv:4:15
	parameter DATAW = 4;
	// Trace: src/VX_stream_xbar.sv:5:15
	parameter ARBITER = "R";
	// Trace: src/VX_stream_xbar.sv:6:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_xbar.sv:7:15
	parameter MAX_FANOUT = 8;
	// Trace: src/VX_stream_xbar.sv:8:15
	parameter PERF_CTR_BITS = $clog2(NUM_INPUTS + 1);
	// Trace: src/VX_stream_xbar.sv:9:15
	parameter IN_WIDTH = (NUM_INPUTS > 1 ? $clog2(NUM_INPUTS) : 1);
	// Trace: src/VX_stream_xbar.sv:10:15
	parameter OUT_WIDTH = (NUM_OUTPUTS > 1 ? $clog2(NUM_OUTPUTS) : 1);
	// Trace: src/VX_stream_xbar.sv:12:5
	input wire clk;
	// Trace: src/VX_stream_xbar.sv:13:5
	input wire reset;
	// Trace: src/VX_stream_xbar.sv:14:5
	input wire [NUM_INPUTS - 1:0] valid_in;
	// Trace: src/VX_stream_xbar.sv:15:5
	input wire [(NUM_INPUTS * DATAW) - 1:0] data_in;
	// Trace: src/VX_stream_xbar.sv:16:5
	input wire [(NUM_INPUTS * OUT_WIDTH) - 1:0] sel_in;
	// Trace: src/VX_stream_xbar.sv:17:5
	output wire [NUM_INPUTS - 1:0] ready_in;
	// Trace: src/VX_stream_xbar.sv:18:5
	output wire [NUM_OUTPUTS - 1:0] valid_out;
	// Trace: src/VX_stream_xbar.sv:19:5
	output wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out;
	// Trace: src/VX_stream_xbar.sv:20:5
	output wire [(NUM_OUTPUTS * IN_WIDTH) - 1:0] sel_out;
	// Trace: src/VX_stream_xbar.sv:21:5
	input wire [NUM_OUTPUTS - 1:0] ready_out;
	// Trace: src/VX_stream_xbar.sv:22:5
	output wire [PERF_CTR_BITS - 1:0] collisions;
	// Trace: src/VX_stream_xbar.sv:24:5
	generate
		if (NUM_INPUTS != 1) begin : g_multi_inputs
			if (NUM_OUTPUTS != 1) begin : g_multiple_outputs
				// Trace: src/VX_stream_xbar.sv:26:13
				wire [(NUM_INPUTS * NUM_OUTPUTS) - 1:0] per_output_valid_in;
				// Trace: src/VX_stream_xbar.sv:27:13
				wire [(NUM_OUTPUTS * NUM_INPUTS) - 1:0] per_output_valid_in_w;
				// Trace: src/VX_stream_xbar.sv:28:13
				wire [(NUM_OUTPUTS * NUM_INPUTS) - 1:0] per_output_ready_in;
				// Trace: src/VX_stream_xbar.sv:29:13
				wire [(NUM_INPUTS * NUM_OUTPUTS) - 1:0] per_output_ready_in_w;
				// Trace: src/VX_stream_xbar.sv:30:13
				VX_transpose #(
					.N(NUM_OUTPUTS),
					.M(NUM_INPUTS)
				) rdy_in_transpose(
					.data_in(per_output_ready_in),
					.data_out(per_output_ready_in_w)
				);
				genvar _gv_i_68;
				for (_gv_i_68 = 0; _gv_i_68 < NUM_INPUTS; _gv_i_68 = _gv_i_68 + 1) begin : g_ready_in
					localparam i = _gv_i_68;
					// Trace: src/VX_stream_xbar.sv:38:17
					assign ready_in[i] = |per_output_ready_in_w[i * NUM_OUTPUTS+:NUM_OUTPUTS];
				end
				genvar _gv_i_69;
				for (_gv_i_69 = 0; _gv_i_69 < NUM_INPUTS; _gv_i_69 = _gv_i_69 + 1) begin : g_sel_in_demux
					localparam i = _gv_i_69;
					// Trace: src/VX_stream_xbar.sv:41:17
					VX_demux #(
						.DATAW(1),
						.N(NUM_OUTPUTS)
					) sel_in_demux(
						.sel_in(sel_in[i * OUT_WIDTH+:OUT_WIDTH]),
						.data_in(valid_in[i]),
						.data_out(per_output_valid_in[i * NUM_OUTPUTS+:NUM_OUTPUTS])
					);
				end
				// Trace: src/VX_stream_xbar.sv:50:13
				VX_transpose #(
					.N(NUM_INPUTS),
					.M(NUM_OUTPUTS)
				) val_in_transpose(
					.data_in(per_output_valid_in),
					.data_out(per_output_valid_in_w)
				);
				genvar _gv_i_70;
				for (_gv_i_70 = 0; _gv_i_70 < NUM_OUTPUTS; _gv_i_70 = _gv_i_70 + 1) begin : g_xbar_arbs
					localparam i = _gv_i_70;
					// Trace: src/VX_stream_xbar.sv:58:17
					VX_stream_arb #(
						.NUM_INPUTS(NUM_INPUTS),
						.NUM_OUTPUTS(1),
						.DATAW(DATAW),
						.ARBITER(ARBITER),
						.MAX_FANOUT(MAX_FANOUT),
						.OUT_BUF(OUT_BUF)
					) xbar_arb(
						.clk(clk),
						.reset(reset),
						.valid_in(per_output_valid_in_w[i * NUM_INPUTS+:NUM_INPUTS]),
						.data_in(data_in),
						.ready_in(per_output_ready_in[i * NUM_INPUTS+:NUM_INPUTS]),
						.valid_out(valid_out[i]),
						.data_out(data_out[i * DATAW+:DATAW]),
						.sel_out(sel_out[i * IN_WIDTH+:IN_WIDTH]),
						.ready_out(ready_out[i])
					);
				end
			end
			else begin : g_one_output
				// Trace: src/VX_stream_xbar.sv:78:13
				VX_stream_arb #(
					.NUM_INPUTS(NUM_INPUTS),
					.NUM_OUTPUTS(1),
					.DATAW(DATAW),
					.ARBITER(ARBITER),
					.MAX_FANOUT(MAX_FANOUT),
					.OUT_BUF(OUT_BUF)
				) xbar_arb(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_in),
					.data_in(data_in),
					.ready_in(ready_in),
					.valid_out(valid_out),
					.data_out(data_out),
					.sel_out(sel_out),
					.ready_out(ready_out)
				);
			end
		end
		else if (NUM_OUTPUTS != 1) begin : g_single_input
			// Trace: src/VX_stream_xbar.sv:98:9
			wire [NUM_OUTPUTS - 1:0] valid_out_w;
			wire [NUM_OUTPUTS - 1:0] ready_out_w;
			// Trace: src/VX_stream_xbar.sv:99:9
			wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out_w;
			// Trace: src/VX_stream_xbar.sv:100:9
			VX_demux #(
				.DATAW(1),
				.N(NUM_OUTPUTS)
			) sel_in_demux(
				.sel_in(sel_in[0+:OUT_WIDTH]),
				.data_in(valid_in[0]),
				.data_out(valid_out_w)
			);
			// Trace: src/VX_stream_xbar.sv:108:9
			assign ready_in[0] = ready_out_w[sel_in[0+:OUT_WIDTH]];
			// Trace: src/VX_stream_xbar.sv:109:9
			assign data_out_w = {NUM_OUTPUTS {data_in[0+:DATAW]}};
			genvar _gv_i_71;
			for (_gv_i_71 = 0; _gv_i_71 < NUM_OUTPUTS; _gv_i_71 = _gv_i_71 + 1) begin : g_out_buf
				localparam i = _gv_i_71;
				// Trace: src/VX_stream_xbar.sv:111:13
				VX_elastic_buffer #(
					.DATAW(DATAW),
					.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
					.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
					.LUTRAM((OUT_BUF & 8) != 0)
				) out_buf(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_out_w[i]),
					.ready_in(ready_out_w[i]),
					.data_in(data_out_w[i * DATAW+:DATAW]),
					.data_out(data_out[i * DATAW+:DATAW]),
					.valid_out(valid_out[i]),
					.ready_out(ready_out[i])
				);
			end
			// Trace: src/VX_stream_xbar.sv:127:9
			assign sel_out = 0;
		end
		else begin : g_passthru
			// Trace: src/VX_stream_xbar.sv:129:9
			VX_elastic_buffer #(
				.DATAW(DATAW),
				.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
				.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
				.LUTRAM((OUT_BUF & 8) != 0)
			) out_buf(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_in),
				.ready_in(ready_in),
				.data_in(data_in),
				.data_out(data_out),
				.valid_out(valid_out),
				.ready_out(ready_out)
			);
			// Trace: src/VX_stream_xbar.sv:144:9
			assign sel_out = 0;
		end
	endgenerate
	// Trace: src/VX_stream_xbar.sv:146:5
	reg [NUM_INPUTS - 1:0] per_cycle_collision;
	reg [NUM_INPUTS - 1:0] per_cycle_collision_r;
	// Trace: src/VX_stream_xbar.sv:147:5
	wire [$clog2(NUM_INPUTS + 1) - 1:0] collision_count;
	// Trace: src/VX_stream_xbar.sv:148:5
	reg [PERF_CTR_BITS - 1:0] collisions_r;
	// Trace: src/VX_stream_xbar.sv:149:5
	always @(*) begin
		// Trace: src/VX_stream_xbar.sv:150:9
		per_cycle_collision = 0;
		// Trace: src/VX_stream_xbar.sv:151:9
		begin : sv2v_autoblock_1
			// Trace: src/VX_stream_xbar.sv:151:14
			integer i;
			// Trace: src/VX_stream_xbar.sv:151:14
			for (i = 0; i < NUM_INPUTS; i = i + 1)
				begin
					// Trace: src/VX_stream_xbar.sv:152:13
					begin : sv2v_autoblock_2
						// Trace: src/VX_stream_xbar.sv:152:18
						integer j;
						// Trace: src/VX_stream_xbar.sv:152:18
						for (j = 1; j < (NUM_INPUTS - i); j = j + 1)
							begin
								// Trace: src/VX_stream_xbar.sv:153:17
								per_cycle_collision[i] = per_cycle_collision[i] | (((valid_in[i] && valid_in[j + i]) && (sel_in[i * OUT_WIDTH+:OUT_WIDTH] == sel_in[(j + i) * OUT_WIDTH+:OUT_WIDTH])) && (ready_in[i] | ready_in[j + i]));
							end
					end
				end
		end
	end
	// Trace: src/VX_stream_xbar.sv:160:5
	// rewrote reg-to-output bindings
	wire [NUM_INPUTS:1] sv2v_tmp___per_cycle_collision_r___data_out;
	always @(*) per_cycle_collision_r = sv2v_tmp___per_cycle_collision_r___data_out;
	VX_pipe_register #(
		.DATAW(NUM_INPUTS),
		.RESETW(0),
		.DEPTH(1)
	) __per_cycle_collision_r__(
		.clk(clk),
		.reset(reset),
		.enable(1'b1),
		.data_in(per_cycle_collision),
		.data_out(sv2v_tmp___per_cycle_collision_r___data_out)
	);
	// Trace: src/VX_stream_xbar.sv:171:5
	VX_popcount #(
		.N(NUM_INPUTS),
		.MODEL(1)
	) __collision_count__(
		.data_in(per_cycle_collision_r),
		.data_out(collision_count)
	);
	// Trace: src/VX_stream_xbar.sv:178:5
	function automatic [PERF_CTR_BITS - 1:0] sv2v_cast_8BEE5;
		input reg [PERF_CTR_BITS - 1:0] inp;
		sv2v_cast_8BEE5 = inp;
	endfunction
	always @(posedge clk)
		// Trace: src/VX_stream_xbar.sv:179:9
		if (reset)
			// Trace: src/VX_stream_xbar.sv:180:13
			collisions_r <= 1'sb0;
		else
			// Trace: src/VX_stream_xbar.sv:182:13
			collisions_r <= collisions_r + sv2v_cast_8BEE5(collision_count);
	// Trace: src/VX_stream_xbar.sv:185:5
	assign collisions = collisions_r;
endmodule
// removed interface: VX_sfu_perf_if
// removed interface: VX_operands_if
// removed module with interface ports: VX_local_mem
module VX_priority_arbiter (
	requests,
	grant_index,
	grant_onehot,
	grant_valid
);
	// Trace: src/VX_priority_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_priority_arbiter.sv:3:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_priority_arbiter.sv:5:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_priority_arbiter.sv:6:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_priority_arbiter.sv:7:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_priority_arbiter.sv:8:5
	output wire grant_valid;
	// Trace: src/VX_priority_arbiter.sv:10:5
	generate
		if (NUM_REQS == 1) begin : g_passthru
			// Trace: src/VX_priority_arbiter.sv:11:9
			assign grant_index = 1'sb0;
			// Trace: src/VX_priority_arbiter.sv:12:9
			assign grant_onehot = requests;
			// Trace: src/VX_priority_arbiter.sv:13:9
			assign grant_valid = requests[0];
		end
		else begin : g_encoder
			// Trace: src/VX_priority_arbiter.sv:15:9
			VX_priority_encoder #(.N(NUM_REQS)) priority_encoder(
				.data_in(requests),
				.index_out(grant_index),
				.onehot_out(grant_onehot),
				.valid_out(grant_valid)
			);
		end
	endgenerate
endmodule
module VX_shift_register (
	clk,
	reset,
	enable,
	data_in,
	data_out
);
	// Trace: src/VX_shift_register.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_shift_register.sv:3:15
	parameter RESETW = 0;
	// Trace: src/VX_shift_register.sv:4:15
	parameter DEPTH = 1;
	// Trace: src/VX_shift_register.sv:5:15
	parameter NUM_TAPS = 1;
	// Trace: src/VX_shift_register.sv:6:15
	parameter TAP_START = 0;
	// Trace: src/VX_shift_register.sv:7:15
	parameter TAP_STRIDE = 1;
	// Trace: src/VX_shift_register.sv:9:5
	input wire clk;
	// Trace: src/VX_shift_register.sv:10:5
	input wire reset;
	// Trace: src/VX_shift_register.sv:11:5
	input wire enable;
	// Trace: src/VX_shift_register.sv:12:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_shift_register.sv:13:5
	output wire [(NUM_TAPS * DATAW) - 1:0] data_out;
	// Trace: src/VX_shift_register.sv:15:5
	generate
		if (DEPTH != 0) begin : g_shift_register
			// Trace: src/VX_shift_register.sv:16:9
			reg [(DEPTH * DATAW) - 1:0] entries;
			// Trace: src/VX_shift_register.sv:17:9
			always @(posedge clk)
				// Trace: src/VX_shift_register.sv:18:13
				begin : sv2v_autoblock_1
					// Trace: src/VX_shift_register.sv:18:18
					integer i;
					// Trace: src/VX_shift_register.sv:18:18
					for (i = 0; i < DATAW; i = i + 1)
						begin
							// Trace: src/VX_shift_register.sv:19:17
							if ((i >= (DATAW - RESETW)) && reset)
								// Trace: src/VX_shift_register.sv:20:21
								begin : sv2v_autoblock_2
									// Trace: src/VX_shift_register.sv:20:26
									integer j;
									// Trace: src/VX_shift_register.sv:20:26
									for (j = 0; j < DEPTH; j = j + 1)
										begin
											// Trace: src/VX_shift_register.sv:21:25
											entries[(j * DATAW) + i] <= 0;
										end
								end
							else if (enable) begin
								// Trace: src/VX_shift_register.sv:23:21
								begin : sv2v_autoblock_3
									// Trace: src/VX_shift_register.sv:23:26
									integer j;
									// Trace: src/VX_shift_register.sv:23:26
									for (j = 1; j < DEPTH; j = j + 1)
										begin
											// Trace: src/VX_shift_register.sv:24:25
											entries[((j - 1) * DATAW) + i] <= entries[(j * DATAW) + i];
										end
								end
								// Trace: src/VX_shift_register.sv:25:21
								entries[((DEPTH - 1) * DATAW) + i] <= data_in[i];
							end
						end
				end
			genvar _gv_i_79;
			for (_gv_i_79 = 0; _gv_i_79 < NUM_TAPS; _gv_i_79 = _gv_i_79 + 1) begin : g_data_out
				localparam i = _gv_i_79;
				// Trace: src/VX_shift_register.sv:30:13
				assign data_out[i * DATAW+:DATAW] = entries[((i * TAP_STRIDE) + TAP_START) * DATAW+:DATAW];
			end
		end
		else begin : g_passthru
			// Trace: src/VX_shift_register.sv:33:9
			assign data_out = data_in;
		end
	endgenerate
endmodule
// removed interface: VX_branch_ctl_if
// removed module with interface ports: VX_mem_arb
// removed module with interface ports: VX_decode
// removed interface: VX_gbar_bus_if
module VX_ipdom_stack (
	clk,
	reset,
	q0,
	q1,
	d,
	d_set,
	q_ptr,
	push,
	pop,
	empty,
	full
);
	// Trace: src/VX_ipdom_stack.sv:2:15
	parameter WIDTH = 1;
	// Trace: src/VX_ipdom_stack.sv:3:15
	parameter DEPTH = 1;
	// Trace: src/VX_ipdom_stack.sv:4:15
	parameter ADDRW = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: src/VX_ipdom_stack.sv:6:5
	input wire clk;
	// Trace: src/VX_ipdom_stack.sv:7:5
	input wire reset;
	// Trace: src/VX_ipdom_stack.sv:8:5
	input wire [WIDTH - 1:0] q0;
	// Trace: src/VX_ipdom_stack.sv:9:5
	input wire [WIDTH - 1:0] q1;
	// Trace: src/VX_ipdom_stack.sv:10:5
	output wire [WIDTH - 1:0] d;
	// Trace: src/VX_ipdom_stack.sv:11:5
	output wire d_set;
	// Trace: src/VX_ipdom_stack.sv:12:5
	output wire [ADDRW - 1:0] q_ptr;
	// Trace: src/VX_ipdom_stack.sv:13:5
	input wire push;
	// Trace: src/VX_ipdom_stack.sv:14:5
	input wire pop;
	// Trace: src/VX_ipdom_stack.sv:15:5
	output wire empty;
	// Trace: src/VX_ipdom_stack.sv:16:5
	output wire full;
	// Trace: src/VX_ipdom_stack.sv:18:5
	reg [ADDRW - 1:0] rd_ptr;
	reg [ADDRW - 1:0] rd_ptr_n;
	reg [ADDRW - 1:0] wr_ptr;
	// Trace: src/VX_ipdom_stack.sv:19:5
	reg empty_r;
	reg full_r;
	// Trace: src/VX_ipdom_stack.sv:20:5
	wire [WIDTH - 1:0] d0;
	wire [WIDTH - 1:0] d1;
	// Trace: src/VX_ipdom_stack.sv:21:5
	wire d_set_r;
	// Trace: src/VX_ipdom_stack.sv:22:5
	function automatic [ADDRW - 1:0] sv2v_cast_8BB5D;
		input reg [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D = inp;
	endfunction
	always @(*) begin
		// Trace: src/VX_ipdom_stack.sv:23:9
		rd_ptr_n = rd_ptr;
		// Trace: src/VX_ipdom_stack.sv:24:9
		if (push)
			// Trace: src/VX_ipdom_stack.sv:25:13
			rd_ptr_n = wr_ptr;
		else if (pop)
			// Trace: src/VX_ipdom_stack.sv:27:13
			rd_ptr_n = rd_ptr - sv2v_cast_8BB5D(d_set_r);
	end
	// Trace: src/VX_ipdom_stack.sv:30:5
	function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
		input reg signed [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D_signed = inp;
	endfunction
	always @(posedge clk)
		// Trace: src/VX_ipdom_stack.sv:31:9
		if (reset) begin
			// Trace: src/VX_ipdom_stack.sv:32:13
			wr_ptr <= 1'sb0;
			// Trace: src/VX_ipdom_stack.sv:33:13
			empty_r <= 1;
			// Trace: src/VX_ipdom_stack.sv:34:13
			full_r <= 0;
			// Trace: src/VX_ipdom_stack.sv:35:13
			rd_ptr <= 1'sb0;
		end
		else begin
			// Trace: src/VX_ipdom_stack.sv:37:13
			if (push) begin
				// Trace: src/VX_ipdom_stack.sv:41:17
				wr_ptr <= wr_ptr + sv2v_cast_8BB5D_signed(1);
				// Trace: src/VX_ipdom_stack.sv:42:17
				empty_r <= 0;
				// Trace: src/VX_ipdom_stack.sv:43:17
				full_r <= sv2v_cast_8BB5D_signed(DEPTH - 1) == wr_ptr;
			end
			else if (pop) begin
				// Trace: src/VX_ipdom_stack.sv:45:17
				wr_ptr <= wr_ptr - sv2v_cast_8BB5D(d_set_r);
				// Trace: src/VX_ipdom_stack.sv:46:17
				empty_r <= (rd_ptr == 0) && d_set_r;
				// Trace: src/VX_ipdom_stack.sv:47:17
				full_r <= 0;
			end
			// Trace: src/VX_ipdom_stack.sv:49:13
			rd_ptr <= rd_ptr_n;
		end
	// Trace: src/VX_ipdom_stack.sv:52:5
	wire [WIDTH * 2:0] qout = (push ? {1'b0, q1, q0} : {1'b1, d1, d0});
	// Trace: src/VX_ipdom_stack.sv:53:5
	VX_dp_ram #(
		.DATAW(1 + (WIDTH * 2)),
		.SIZE(DEPTH),
		.OUT_REG(1),
		.RDW_MODE("R")
	) ipdom_store(
		.clk(clk),
		.reset(reset),
		.read(1'b1),
		.write(push || pop),
		.wren(1'b1),
		.waddr((push ? wr_ptr : rd_ptr)),
		.wdata(qout),
		.raddr(rd_ptr_n),
		.rdata({d_set_r, d1, d0})
	);
	// Trace: src/VX_ipdom_stack.sv:69:5
	assign d = (d_set_r ? d0 : d1);
	// Trace: src/VX_ipdom_stack.sv:70:5
	assign d_set = ~d_set_r;
	// Trace: src/VX_ipdom_stack.sv:71:5
	assign q_ptr = wr_ptr;
	// Trace: src/VX_ipdom_stack.sv:72:5
	assign empty = empty_r;
	// Trace: src/VX_ipdom_stack.sv:73:5
	assign full = full_r;
endmodule
// removed interface: VX_commit_sched_if
module VX_multiplier (
	clk,
	enable,
	dataa,
	datab,
	result
);
	// Trace: src/VX_multiplier.sv:2:15
	parameter A_WIDTH = 1;
	// Trace: src/VX_multiplier.sv:3:15
	parameter B_WIDTH = A_WIDTH;
	// Trace: src/VX_multiplier.sv:4:15
	parameter R_WIDTH = A_WIDTH + B_WIDTH;
	// Trace: src/VX_multiplier.sv:5:15
	parameter SIGNED = 0;
	// Trace: src/VX_multiplier.sv:6:15
	parameter LATENCY = 0;
	// Trace: src/VX_multiplier.sv:8:5
	input wire clk;
	// Trace: src/VX_multiplier.sv:9:5
	input wire enable;
	// Trace: src/VX_multiplier.sv:10:5
	input wire [A_WIDTH - 1:0] dataa;
	// Trace: src/VX_multiplier.sv:11:5
	input wire [B_WIDTH - 1:0] datab;
	// Trace: src/VX_multiplier.sv:12:5
	output wire [R_WIDTH - 1:0] result;
	// Trace: src/VX_multiplier.sv:14:5
	wire [R_WIDTH - 1:0] prod_w;
	// Trace: src/VX_multiplier.sv:15:5
	function automatic [R_WIDTH - 1:0] sv2v_cast_875D6;
		input reg [R_WIDTH - 1:0] inp;
		sv2v_cast_875D6 = inp;
	endfunction
	function automatic signed [R_WIDTH - 1:0] sv2v_cast_875D6_signed;
		input reg signed [R_WIDTH - 1:0] inp;
		sv2v_cast_875D6_signed = inp;
	endfunction
	generate
		if (SIGNED != 0) begin : g_prod_s
			// Trace: src/VX_multiplier.sv:16:9
			assign prod_w = sv2v_cast_875D6_signed($signed(dataa) * $signed(datab));
		end
		else begin : g_prod_u
			// Trace: src/VX_multiplier.sv:18:9
			assign prod_w = sv2v_cast_875D6(dataa * datab);
		end
	endgenerate
	// Trace: src/VX_multiplier.sv:20:5
	generate
		if (LATENCY == 0) begin : g_passthru
			// Trace: src/VX_multiplier.sv:21:9
			assign result = prod_w;
		end
		else begin : g_latency
			// Trace: src/VX_multiplier.sv:23:9
			reg [(LATENCY * R_WIDTH) - 1:0] prod_r;
			// Trace: src/VX_multiplier.sv:24:9
			always @(posedge clk)
				// Trace: src/VX_multiplier.sv:25:13
				if (enable) begin
					// Trace: src/VX_multiplier.sv:26:17
					prod_r[0+:R_WIDTH] <= prod_w;
					// Trace: src/VX_multiplier.sv:27:17
					begin : sv2v_autoblock_1
						// Trace: src/VX_multiplier.sv:27:22
						integer i;
						// Trace: src/VX_multiplier.sv:27:22
						for (i = 1; i < LATENCY; i = i + 1)
							begin
								// Trace: src/VX_multiplier.sv:28:21
								prod_r[i * R_WIDTH+:R_WIDTH] <= prod_r[(i - 1) * R_WIDTH+:R_WIDTH];
							end
					end
				end
			// Trace: src/VX_multiplier.sv:32:9
			assign result = prod_r[(LATENCY - 1) * R_WIDTH+:R_WIDTH];
		end
	endgenerate
endmodule
// removed module with interface ports: VX_lsu_mem_arb
// removed module with interface ports: VX_core
module VX_bits_insert (
	data_in,
	ins_in,
	data_out
);
	// Trace: src/VX_bits_insert.sv:2:15
	parameter N = 1;
	// Trace: src/VX_bits_insert.sv:3:15
	parameter S = 1;
	// Trace: src/VX_bits_insert.sv:4:15
	parameter POS = 0;
	// Trace: src/VX_bits_insert.sv:6:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_bits_insert.sv:7:5
	input wire [(S > 0 ? S : 1) - 1:0] ins_in;
	// Trace: src/VX_bits_insert.sv:8:5
	output wire [(N + S) - 1:0] data_out;
	// Trace: src/VX_bits_insert.sv:10:5
	generate
		if (S == 0) begin : g_passthru
			// Trace: src/VX_bits_insert.sv:11:9
			assign data_out = data_in;
		end
		else begin : g_insert
			if (POS == 0) begin : g_pos_0
				// Trace: src/VX_bits_insert.sv:14:13
				assign data_out = {data_in, ins_in};
			end
			else if (POS == N) begin : g_pos_N
				// Trace: src/VX_bits_insert.sv:16:13
				assign data_out = {ins_in, data_in};
			end
			else begin : g_pos
				// Trace: src/VX_bits_insert.sv:18:13
				assign data_out = {data_in[N - 1:POS], ins_in, data_in[POS - 1:0]};
			end
		end
	endgenerate
endmodule
module VX_mem_scheduler (
	clk,
	reset,
	core_req_valid,
	core_req_rw,
	core_req_mask,
	core_req_byteen,
	core_req_addr,
	core_req_flags,
	core_req_data,
	core_req_tag,
	core_req_ready,
	core_req_empty,
	core_req_wr_notify,
	core_rsp_valid,
	core_rsp_mask,
	core_rsp_data,
	core_rsp_tag,
	core_rsp_sop,
	core_rsp_eop,
	core_rsp_ready,
	mem_req_valid,
	mem_req_rw,
	mem_req_mask,
	mem_req_byteen,
	mem_req_addr,
	mem_req_flags,
	mem_req_data,
	mem_req_tag,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_mask,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready
);
	// Trace: src/VX_mem_scheduler.sv:2:15
	parameter INSTANCE_ID = "";
	// Trace: src/VX_mem_scheduler.sv:3:15
	parameter CORE_REQS = 1;
	// Trace: src/VX_mem_scheduler.sv:4:15
	parameter MEM_CHANNELS = 1;
	// Trace: src/VX_mem_scheduler.sv:5:15
	parameter WORD_SIZE = 4;
	// Trace: src/VX_mem_scheduler.sv:6:15
	parameter LINE_SIZE = WORD_SIZE;
	// Trace: src/VX_mem_scheduler.sv:7:15
	parameter ADDR_WIDTH = 32 - $clog2(WORD_SIZE);
	// Trace: src/VX_mem_scheduler.sv:8:15
	parameter FLAGS_WIDTH = 0;
	// Trace: src/VX_mem_scheduler.sv:9:15
	parameter TAG_WIDTH = 8;
	// Trace: src/VX_mem_scheduler.sv:10:15
	parameter UUID_WIDTH = 0;
	// Trace: src/VX_mem_scheduler.sv:11:15
	parameter CORE_QUEUE_SIZE = 8;
	// Trace: src/VX_mem_scheduler.sv:12:15
	parameter MEM_QUEUE_SIZE = CORE_QUEUE_SIZE;
	// Trace: src/VX_mem_scheduler.sv:13:15
	parameter RSP_PARTIAL = 0;
	// Trace: src/VX_mem_scheduler.sv:14:15
	parameter CORE_OUT_BUF = 0;
	// Trace: src/VX_mem_scheduler.sv:15:15
	parameter MEM_OUT_BUF = 0;
	// Trace: src/VX_mem_scheduler.sv:16:15
	parameter WORD_WIDTH = WORD_SIZE * 8;
	// Trace: src/VX_mem_scheduler.sv:17:15
	parameter LINE_WIDTH = LINE_SIZE * 8;
	// Trace: src/VX_mem_scheduler.sv:18:15
	parameter COALESCE_ENABLE = (CORE_REQS > 1) && (LINE_SIZE != WORD_SIZE);
	// Trace: src/VX_mem_scheduler.sv:19:15
	parameter PER_LINE_REQS = LINE_SIZE / WORD_SIZE;
	// Trace: src/VX_mem_scheduler.sv:20:15
	parameter MERGED_REQS = CORE_REQS / PER_LINE_REQS;
	// Trace: src/VX_mem_scheduler.sv:21:15
	parameter MEM_BATCHES = ((MERGED_REQS + MEM_CHANNELS) - 1) / MEM_CHANNELS;
	// Trace: src/VX_mem_scheduler.sv:22:15
	parameter MEM_BATCH_BITS = $clog2(MEM_BATCHES);
	// Trace: src/VX_mem_scheduler.sv:23:15
	parameter MEM_QUEUE_ADDRW = $clog2((COALESCE_ENABLE ? MEM_QUEUE_SIZE : CORE_QUEUE_SIZE));
	// Trace: src/VX_mem_scheduler.sv:24:15
	parameter MEM_ADDR_WIDTH = ADDR_WIDTH - $clog2(PER_LINE_REQS);
	// Trace: src/VX_mem_scheduler.sv:25:15
	parameter MEM_TAG_WIDTH = (UUID_WIDTH + MEM_QUEUE_ADDRW) + MEM_BATCH_BITS;
	// Trace: src/VX_mem_scheduler.sv:27:5
	input wire clk;
	// Trace: src/VX_mem_scheduler.sv:28:5
	input wire reset;
	// Trace: src/VX_mem_scheduler.sv:29:5
	input wire core_req_valid;
	// Trace: src/VX_mem_scheduler.sv:30:5
	input wire core_req_rw;
	// Trace: src/VX_mem_scheduler.sv:31:5
	input wire [CORE_REQS - 1:0] core_req_mask;
	// Trace: src/VX_mem_scheduler.sv:32:5
	input wire [(CORE_REQS * WORD_SIZE) - 1:0] core_req_byteen;
	// Trace: src/VX_mem_scheduler.sv:33:5
	input wire [(CORE_REQS * ADDR_WIDTH) - 1:0] core_req_addr;
	// Trace: src/VX_mem_scheduler.sv:34:5
	input wire [(CORE_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] core_req_flags;
	// Trace: src/VX_mem_scheduler.sv:35:5
	input wire [(CORE_REQS * WORD_WIDTH) - 1:0] core_req_data;
	// Trace: src/VX_mem_scheduler.sv:36:5
	input wire [TAG_WIDTH - 1:0] core_req_tag;
	// Trace: src/VX_mem_scheduler.sv:37:5
	output wire core_req_ready;
	// Trace: src/VX_mem_scheduler.sv:38:5
	output wire core_req_empty;
	// Trace: src/VX_mem_scheduler.sv:39:5
	output wire core_req_wr_notify;
	// Trace: src/VX_mem_scheduler.sv:40:5
	output wire core_rsp_valid;
	// Trace: src/VX_mem_scheduler.sv:41:5
	output wire [CORE_REQS - 1:0] core_rsp_mask;
	// Trace: src/VX_mem_scheduler.sv:42:5
	output wire [(CORE_REQS * WORD_WIDTH) - 1:0] core_rsp_data;
	// Trace: src/VX_mem_scheduler.sv:43:5
	output wire [TAG_WIDTH - 1:0] core_rsp_tag;
	// Trace: src/VX_mem_scheduler.sv:44:5
	output wire core_rsp_sop;
	// Trace: src/VX_mem_scheduler.sv:45:5
	output wire core_rsp_eop;
	// Trace: src/VX_mem_scheduler.sv:46:5
	input wire core_rsp_ready;
	// Trace: src/VX_mem_scheduler.sv:47:5
	output wire mem_req_valid;
	// Trace: src/VX_mem_scheduler.sv:48:5
	output wire mem_req_rw;
	// Trace: src/VX_mem_scheduler.sv:49:5
	output wire [MEM_CHANNELS - 1:0] mem_req_mask;
	// Trace: src/VX_mem_scheduler.sv:50:5
	output wire [(MEM_CHANNELS * LINE_SIZE) - 1:0] mem_req_byteen;
	// Trace: src/VX_mem_scheduler.sv:51:5
	output wire [(MEM_CHANNELS * MEM_ADDR_WIDTH) - 1:0] mem_req_addr;
	// Trace: src/VX_mem_scheduler.sv:52:5
	output wire [(MEM_CHANNELS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] mem_req_flags;
	// Trace: src/VX_mem_scheduler.sv:53:5
	output wire [(MEM_CHANNELS * LINE_WIDTH) - 1:0] mem_req_data;
	// Trace: src/VX_mem_scheduler.sv:54:5
	output wire [MEM_TAG_WIDTH - 1:0] mem_req_tag;
	// Trace: src/VX_mem_scheduler.sv:55:5
	input wire mem_req_ready;
	// Trace: src/VX_mem_scheduler.sv:56:5
	input wire mem_rsp_valid;
	// Trace: src/VX_mem_scheduler.sv:57:5
	input wire [MEM_CHANNELS - 1:0] mem_rsp_mask;
	// Trace: src/VX_mem_scheduler.sv:58:5
	input wire [(MEM_CHANNELS * LINE_WIDTH) - 1:0] mem_rsp_data;
	// Trace: src/VX_mem_scheduler.sv:59:5
	input wire [MEM_TAG_WIDTH - 1:0] mem_rsp_tag;
	// Trace: src/VX_mem_scheduler.sv:60:5
	output wire mem_rsp_ready;
	// Trace: src/VX_mem_scheduler.sv:62:5
	localparam BATCH_SEL_WIDTH = (MEM_BATCH_BITS > 0 ? MEM_BATCH_BITS : 1);
	// Trace: src/VX_mem_scheduler.sv:63:5
	localparam STALL_TIMEOUT = 10000000;
	// Trace: src/VX_mem_scheduler.sv:64:5
	localparam CORE_QUEUE_ADDRW = $clog2(CORE_QUEUE_SIZE);
	// Trace: src/VX_mem_scheduler.sv:65:5
	localparam TAG_ID_WIDTH = TAG_WIDTH - UUID_WIDTH;
	// Trace: src/VX_mem_scheduler.sv:66:5
	localparam REQQ_TAG_WIDTH = UUID_WIDTH + CORE_QUEUE_ADDRW;
	// Trace: src/VX_mem_scheduler.sv:67:5
	localparam MERGED_TAG_WIDTH = UUID_WIDTH + MEM_QUEUE_ADDRW;
	// Trace: src/VX_mem_scheduler.sv:68:5
	localparam CORE_CHANNELS = (COALESCE_ENABLE ? CORE_REQS : MEM_CHANNELS);
	// Trace: src/VX_mem_scheduler.sv:69:5
	localparam CORE_BATCHES = (COALESCE_ENABLE ? 1 : MEM_BATCHES);
	// Trace: src/VX_mem_scheduler.sv:70:5
	localparam CORE_BATCH_BITS = $clog2(CORE_BATCHES);
	// Trace: src/VX_mem_scheduler.sv:71:5
	wire ibuf_push;
	// Trace: src/VX_mem_scheduler.sv:72:5
	wire ibuf_pop;
	// Trace: src/VX_mem_scheduler.sv:73:5
	wire [CORE_QUEUE_ADDRW - 1:0] ibuf_waddr;
	// Trace: src/VX_mem_scheduler.sv:74:5
	wire [CORE_QUEUE_ADDRW - 1:0] ibuf_raddr;
	// Trace: src/VX_mem_scheduler.sv:75:5
	wire ibuf_full;
	// Trace: src/VX_mem_scheduler.sv:76:5
	wire ibuf_empty;
	// Trace: src/VX_mem_scheduler.sv:77:5
	wire [TAG_ID_WIDTH - 1:0] ibuf_din;
	// Trace: src/VX_mem_scheduler.sv:78:5
	wire [TAG_ID_WIDTH - 1:0] ibuf_dout;
	// Trace: src/VX_mem_scheduler.sv:79:5
	wire reqq_valid;
	// Trace: src/VX_mem_scheduler.sv:80:5
	wire [CORE_REQS - 1:0] reqq_mask;
	// Trace: src/VX_mem_scheduler.sv:81:5
	wire reqq_rw;
	// Trace: src/VX_mem_scheduler.sv:82:5
	wire [(CORE_REQS * WORD_SIZE) - 1:0] reqq_byteen;
	// Trace: src/VX_mem_scheduler.sv:83:5
	wire [(CORE_REQS * ADDR_WIDTH) - 1:0] reqq_addr;
	// Trace: src/VX_mem_scheduler.sv:84:5
	wire [(CORE_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] reqq_flags;
	// Trace: src/VX_mem_scheduler.sv:85:5
	wire [(CORE_REQS * WORD_WIDTH) - 1:0] reqq_data;
	// Trace: src/VX_mem_scheduler.sv:86:5
	wire [REQQ_TAG_WIDTH - 1:0] reqq_tag;
	// Trace: src/VX_mem_scheduler.sv:87:5
	wire reqq_ready;
	// Trace: src/VX_mem_scheduler.sv:88:5
	wire reqq_valid_s;
	// Trace: src/VX_mem_scheduler.sv:89:5
	wire [MERGED_REQS - 1:0] reqq_mask_s;
	// Trace: src/VX_mem_scheduler.sv:90:5
	wire reqq_rw_s;
	// Trace: src/VX_mem_scheduler.sv:91:5
	wire [(MERGED_REQS * LINE_SIZE) - 1:0] reqq_byteen_s;
	// Trace: src/VX_mem_scheduler.sv:92:5
	wire [(MERGED_REQS * MEM_ADDR_WIDTH) - 1:0] reqq_addr_s;
	// Trace: src/VX_mem_scheduler.sv:93:5
	wire [(MERGED_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] reqq_flags_s;
	// Trace: src/VX_mem_scheduler.sv:94:5
	wire [(MERGED_REQS * LINE_WIDTH) - 1:0] reqq_data_s;
	// Trace: src/VX_mem_scheduler.sv:95:5
	wire [MERGED_TAG_WIDTH - 1:0] reqq_tag_s;
	// Trace: src/VX_mem_scheduler.sv:96:5
	wire reqq_ready_s;
	// Trace: src/VX_mem_scheduler.sv:97:5
	wire mem_req_valid_s;
	// Trace: src/VX_mem_scheduler.sv:98:5
	wire [MEM_CHANNELS - 1:0] mem_req_mask_s;
	// Trace: src/VX_mem_scheduler.sv:99:5
	wire mem_req_rw_s;
	// Trace: src/VX_mem_scheduler.sv:100:5
	wire [(MEM_CHANNELS * LINE_SIZE) - 1:0] mem_req_byteen_s;
	// Trace: src/VX_mem_scheduler.sv:101:5
	wire [(MEM_CHANNELS * MEM_ADDR_WIDTH) - 1:0] mem_req_addr_s;
	// Trace: src/VX_mem_scheduler.sv:102:5
	wire [(MEM_CHANNELS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] mem_req_flags_s;
	// Trace: src/VX_mem_scheduler.sv:103:5
	wire [(MEM_CHANNELS * LINE_WIDTH) - 1:0] mem_req_data_s;
	// Trace: src/VX_mem_scheduler.sv:104:5
	wire [MEM_TAG_WIDTH - 1:0] mem_req_tag_s;
	// Trace: src/VX_mem_scheduler.sv:105:5
	wire mem_req_ready_s;
	// Trace: src/VX_mem_scheduler.sv:106:5
	wire mem_rsp_valid_s;
	// Trace: src/VX_mem_scheduler.sv:107:5
	wire [CORE_CHANNELS - 1:0] mem_rsp_mask_s;
	// Trace: src/VX_mem_scheduler.sv:108:5
	wire [(CORE_CHANNELS * WORD_WIDTH) - 1:0] mem_rsp_data_s;
	// Trace: src/VX_mem_scheduler.sv:109:5
	wire [MEM_TAG_WIDTH - 1:0] mem_rsp_tag_s;
	// Trace: src/VX_mem_scheduler.sv:110:5
	wire mem_rsp_ready_s;
	// Trace: src/VX_mem_scheduler.sv:111:5
	wire crsp_valid;
	// Trace: src/VX_mem_scheduler.sv:112:5
	wire [CORE_REQS - 1:0] crsp_mask;
	// Trace: src/VX_mem_scheduler.sv:113:5
	wire [(CORE_REQS * WORD_WIDTH) - 1:0] crsp_data;
	// Trace: src/VX_mem_scheduler.sv:114:5
	wire [TAG_WIDTH - 1:0] crsp_tag;
	// Trace: src/VX_mem_scheduler.sv:115:5
	wire crsp_sop;
	// Trace: src/VX_mem_scheduler.sv:116:5
	wire crsp_eop;
	// Trace: src/VX_mem_scheduler.sv:117:5
	wire crsp_ready;
	// Trace: src/VX_mem_scheduler.sv:118:5
	wire req_sent_all;
	// Trace: src/VX_mem_scheduler.sv:119:5
	wire ibuf_ready = core_req_rw || ~ibuf_full;
	// Trace: src/VX_mem_scheduler.sv:120:5
	wire reqq_valid_in = core_req_valid && ibuf_ready;
	// Trace: src/VX_mem_scheduler.sv:121:5
	wire reqq_ready_in;
	// Trace: src/VX_mem_scheduler.sv:122:5
	wire [REQQ_TAG_WIDTH - 1:0] reqq_tag_u;
	// Trace: src/VX_mem_scheduler.sv:123:5
	generate
		if (UUID_WIDTH != 0) begin : g_reqq_tag_u_uuid
			// Trace: src/VX_mem_scheduler.sv:124:9
			assign reqq_tag_u = {core_req_tag[TAG_WIDTH - 1-:UUID_WIDTH], ibuf_waddr};
		end
		else begin : g_reqq_tag_u
			// Trace: src/VX_mem_scheduler.sv:126:9
			assign reqq_tag_u = ibuf_waddr;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:128:5
	VX_elastic_buffer #(
		.DATAW((1 + (CORE_REQS * ((((1 + WORD_SIZE) + ADDR_WIDTH) + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + WORD_WIDTH))) + REQQ_TAG_WIDTH),
		.SIZE(CORE_QUEUE_SIZE),
		.OUT_REG(1)
	) req_queue(
		.clk(clk),
		.reset(reset),
		.valid_in(reqq_valid_in),
		.ready_in(reqq_ready_in),
		.data_in({core_req_rw, core_req_mask, core_req_byteen, core_req_addr, core_req_flags, core_req_data, reqq_tag_u}),
		.data_out({reqq_rw, reqq_mask, reqq_byteen, reqq_addr, reqq_flags, reqq_data, reqq_tag}),
		.valid_out(reqq_valid),
		.ready_out(reqq_ready)
	);
	// Trace: src/VX_mem_scheduler.sv:142:5
	assign core_req_ready = reqq_ready_in && ibuf_ready;
	// Trace: src/VX_mem_scheduler.sv:143:5
	assign core_req_empty = !reqq_valid && ibuf_empty;
	// Trace: src/VX_mem_scheduler.sv:144:5
	assign core_req_wr_notify = (reqq_valid && reqq_ready) && reqq_rw;
	// Trace: src/VX_mem_scheduler.sv:145:5
	wire core_req_fire = core_req_valid && core_req_ready;
	// Trace: src/VX_mem_scheduler.sv:146:5
	wire crsp_fire = crsp_valid && crsp_ready;
	// Trace: src/VX_mem_scheduler.sv:147:5
	assign ibuf_push = core_req_fire && ~core_req_rw;
	// Trace: src/VX_mem_scheduler.sv:148:5
	assign ibuf_pop = crsp_fire && crsp_eop;
	// Trace: src/VX_mem_scheduler.sv:149:5
	assign ibuf_raddr = mem_rsp_tag_s[CORE_BATCH_BITS+:CORE_QUEUE_ADDRW];
	// Trace: src/VX_mem_scheduler.sv:150:5
	assign ibuf_din = core_req_tag[TAG_ID_WIDTH - 1:0];
	// Trace: src/VX_mem_scheduler.sv:151:5
	VX_index_buffer #(
		.DATAW(TAG_ID_WIDTH),
		.SIZE(CORE_QUEUE_SIZE)
	) req_ibuf(
		.clk(clk),
		.reset(reset),
		.acquire_en(ibuf_push),
		.write_addr(ibuf_waddr),
		.write_data(ibuf_din),
		.read_data(ibuf_dout),
		.read_addr(ibuf_raddr),
		.release_en(ibuf_pop),
		.full(ibuf_full),
		.empty(ibuf_empty)
	);
	// Trace: src/VX_mem_scheduler.sv:166:5
	generate
		if (COALESCE_ENABLE) begin : g_coalescer
			// Trace: src/VX_mem_scheduler.sv:167:9
			VX_mem_coalescer #(
				.INSTANCE_ID(""),
				.NUM_REQS(CORE_REQS),
				.DATA_IN_SIZE(WORD_SIZE),
				.DATA_OUT_SIZE(LINE_SIZE),
				.ADDR_WIDTH(ADDR_WIDTH),
				.FLAGS_WIDTH(FLAGS_WIDTH),
				.TAG_WIDTH(REQQ_TAG_WIDTH),
				.UUID_WIDTH(UUID_WIDTH),
				.QUEUE_SIZE(MEM_QUEUE_SIZE)
			) coalescer(
				.clk(clk),
				.reset(reset),
				.in_req_valid(reqq_valid),
				.in_req_mask(reqq_mask),
				.in_req_rw(reqq_rw),
				.in_req_byteen(reqq_byteen),
				.in_req_addr(reqq_addr),
				.in_req_flags(reqq_flags),
				.in_req_data(reqq_data),
				.in_req_tag(reqq_tag),
				.in_req_ready(reqq_ready),
				.in_rsp_valid(mem_rsp_valid_s),
				.in_rsp_mask(mem_rsp_mask_s),
				.in_rsp_data(mem_rsp_data_s),
				.in_rsp_tag(mem_rsp_tag_s),
				.in_rsp_ready(mem_rsp_ready_s),
				.out_req_valid(reqq_valid_s),
				.out_req_mask(reqq_mask_s),
				.out_req_rw(reqq_rw_s),
				.out_req_byteen(reqq_byteen_s),
				.out_req_addr(reqq_addr_s),
				.out_req_flags(reqq_flags_s),
				.out_req_data(reqq_data_s),
				.out_req_tag(reqq_tag_s),
				.out_req_ready(reqq_ready_s),
				.out_rsp_valid(mem_rsp_valid),
				.out_rsp_mask(mem_rsp_mask),
				.out_rsp_data(mem_rsp_data),
				.out_rsp_tag(mem_rsp_tag),
				.out_rsp_ready(mem_rsp_ready)
			);
		end
		else begin : g_no_coalescer
			// Trace: src/VX_mem_scheduler.sv:210:9
			assign reqq_valid_s = reqq_valid;
			// Trace: src/VX_mem_scheduler.sv:211:9
			assign reqq_mask_s = reqq_mask;
			// Trace: src/VX_mem_scheduler.sv:212:9
			assign reqq_rw_s = reqq_rw;
			// Trace: src/VX_mem_scheduler.sv:213:9
			assign reqq_byteen_s = reqq_byteen;
			// Trace: src/VX_mem_scheduler.sv:214:9
			assign reqq_addr_s = reqq_addr;
			// Trace: src/VX_mem_scheduler.sv:215:9
			assign reqq_flags_s = reqq_flags;
			// Trace: src/VX_mem_scheduler.sv:216:9
			assign reqq_data_s = reqq_data;
			// Trace: src/VX_mem_scheduler.sv:217:9
			assign reqq_tag_s = reqq_tag;
			// Trace: src/VX_mem_scheduler.sv:218:9
			assign reqq_ready = reqq_ready_s;
			// Trace: src/VX_mem_scheduler.sv:219:9
			assign mem_rsp_valid_s = mem_rsp_valid;
			// Trace: src/VX_mem_scheduler.sv:220:9
			assign mem_rsp_mask_s = mem_rsp_mask;
			// Trace: src/VX_mem_scheduler.sv:221:9
			assign mem_rsp_data_s = mem_rsp_data;
			// Trace: src/VX_mem_scheduler.sv:222:9
			assign mem_rsp_tag_s = mem_rsp_tag;
			// Trace: src/VX_mem_scheduler.sv:223:9
			assign mem_rsp_ready = mem_rsp_ready_s;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:225:5
	wire [(MEM_BATCHES * MEM_CHANNELS) - 1:0] mem_req_mask_b;
	// Trace: src/VX_mem_scheduler.sv:226:5
	wire [((MEM_BATCHES * MEM_CHANNELS) * LINE_SIZE) - 1:0] mem_req_byteen_b;
	// Trace: src/VX_mem_scheduler.sv:227:5
	wire [((MEM_BATCHES * MEM_CHANNELS) * MEM_ADDR_WIDTH) - 1:0] mem_req_addr_b;
	// Trace: src/VX_mem_scheduler.sv:228:5
	wire [((MEM_BATCHES * MEM_CHANNELS) * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] mem_req_flags_b;
	// Trace: src/VX_mem_scheduler.sv:229:5
	wire [((MEM_BATCHES * MEM_CHANNELS) * LINE_WIDTH) - 1:0] mem_req_data_b;
	// Trace: src/VX_mem_scheduler.sv:230:5
	wire [BATCH_SEL_WIDTH - 1:0] req_batch_idx;
	// Trace: src/VX_mem_scheduler.sv:231:5
	genvar _gv_i_90;
	generate
		for (_gv_i_90 = 0; _gv_i_90 < MEM_BATCHES; _gv_i_90 = _gv_i_90 + 1) begin : g_mem_req_data_b
			localparam i = _gv_i_90;
			genvar _gv_j_8;
			for (_gv_j_8 = 0; _gv_j_8 < MEM_CHANNELS; _gv_j_8 = _gv_j_8 + 1) begin : g_j
				localparam j = _gv_j_8;
				// Trace: src/VX_mem_scheduler.sv:233:13
				localparam r = (i * MEM_CHANNELS) + j;
				if (r < MERGED_REQS) begin : g_valid
					// Trace: src/VX_mem_scheduler.sv:235:17
					assign mem_req_mask_b[(i * MEM_CHANNELS) + j] = reqq_mask_s[r];
					// Trace: src/VX_mem_scheduler.sv:236:17
					assign mem_req_byteen_b[((i * MEM_CHANNELS) + j) * LINE_SIZE+:LINE_SIZE] = reqq_byteen_s[r * LINE_SIZE+:LINE_SIZE];
					// Trace: src/VX_mem_scheduler.sv:237:17
					assign mem_req_addr_b[((i * MEM_CHANNELS) + j) * MEM_ADDR_WIDTH+:MEM_ADDR_WIDTH] = reqq_addr_s[r * MEM_ADDR_WIDTH+:MEM_ADDR_WIDTH];
					// Trace: src/VX_mem_scheduler.sv:238:17
					assign mem_req_flags_b[((i * MEM_CHANNELS) + j) * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)] = reqq_flags_s[r * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)];
					// Trace: src/VX_mem_scheduler.sv:239:17
					assign mem_req_data_b[((i * MEM_CHANNELS) + j) * LINE_WIDTH+:LINE_WIDTH] = reqq_data_s[r * LINE_WIDTH+:LINE_WIDTH];
				end
				else begin : g_padding
					// Trace: src/VX_mem_scheduler.sv:241:17
					assign mem_req_mask_b[(i * MEM_CHANNELS) + j] = 0;
					// Trace: src/VX_mem_scheduler.sv:242:17
					assign mem_req_byteen_b[((i * MEM_CHANNELS) + j) * LINE_SIZE+:LINE_SIZE] = 1'sb0;
					// Trace: src/VX_mem_scheduler.sv:243:17
					assign mem_req_addr_b[((i * MEM_CHANNELS) + j) * MEM_ADDR_WIDTH+:MEM_ADDR_WIDTH] = 1'sb0;
					// Trace: src/VX_mem_scheduler.sv:244:17
					assign mem_req_flags_b[((i * MEM_CHANNELS) + j) * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)] = 1'sb0;
					// Trace: src/VX_mem_scheduler.sv:245:17
					assign mem_req_data_b[((i * MEM_CHANNELS) + j) * LINE_WIDTH+:LINE_WIDTH] = 1'sb0;
				end
			end
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:249:5
	assign mem_req_mask_s = mem_req_mask_b[req_batch_idx * MEM_CHANNELS+:MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:250:5
	assign mem_req_rw_s = reqq_rw_s;
	// Trace: src/VX_mem_scheduler.sv:251:5
	assign mem_req_byteen_s = mem_req_byteen_b[LINE_SIZE * (req_batch_idx * MEM_CHANNELS)+:LINE_SIZE * MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:252:5
	assign mem_req_addr_s = mem_req_addr_b[MEM_ADDR_WIDTH * (req_batch_idx * MEM_CHANNELS)+:MEM_ADDR_WIDTH * MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:253:5
	assign mem_req_flags_s = mem_req_flags_b[(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) * (req_batch_idx * MEM_CHANNELS)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) * MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:254:5
	assign mem_req_data_s = mem_req_data_b[LINE_WIDTH * (req_batch_idx * MEM_CHANNELS)+:LINE_WIDTH * MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:255:5
	function automatic signed [MEM_BATCH_BITS - 1:0] sv2v_cast_F385D_signed;
		input reg signed [MEM_BATCH_BITS - 1:0] inp;
		sv2v_cast_F385D_signed = inp;
	endfunction
	generate
		if (MEM_BATCHES != 1) begin : g_batch
			// Trace: src/VX_mem_scheduler.sv:256:9
			reg [MEM_BATCH_BITS - 1:0] req_batch_idx_r;
			// Trace: src/VX_mem_scheduler.sv:257:9
			wire is_degenerate_batch = ~(|mem_req_mask_s);
			// Trace: src/VX_mem_scheduler.sv:258:9
			wire mem_req_valid_b = reqq_valid_s && ~is_degenerate_batch;
			// Trace: src/VX_mem_scheduler.sv:259:9
			wire mem_req_ready_b = mem_req_ready_s || is_degenerate_batch;
			// Trace: src/VX_mem_scheduler.sv:260:9
			always @(posedge clk)
				// Trace: src/VX_mem_scheduler.sv:261:13
				if (reset)
					// Trace: src/VX_mem_scheduler.sv:262:17
					req_batch_idx_r <= 1'sb0;
				else
					// Trace: src/VX_mem_scheduler.sv:264:17
					if (reqq_valid_s && mem_req_ready_b) begin
						begin
							// Trace: src/VX_mem_scheduler.sv:265:21
							if (req_sent_all)
								// Trace: src/VX_mem_scheduler.sv:266:25
								req_batch_idx_r <= 1'sb0;
							else
								// Trace: src/VX_mem_scheduler.sv:268:25
								req_batch_idx_r <= req_batch_idx_r + sv2v_cast_F385D_signed(1);
						end
					end
			// Trace: src/VX_mem_scheduler.sv:273:9
			wire [MEM_BATCHES - 1:0] req_batch_valids;
			// Trace: src/VX_mem_scheduler.sv:274:9
			wire [(MEM_BATCHES * MEM_BATCH_BITS) - 1:0] req_batch_idxs;
			// Trace: src/VX_mem_scheduler.sv:275:9
			wire [MEM_BATCH_BITS - 1:0] req_batch_idx_last;
			genvar _gv_i_91;
			for (_gv_i_91 = 0; _gv_i_91 < MEM_BATCHES; _gv_i_91 = _gv_i_91 + 1) begin : g_req_batch
				localparam i = _gv_i_91;
				// Trace: src/VX_mem_scheduler.sv:277:13
				assign req_batch_valids[i] = |mem_req_mask_b[i * MEM_CHANNELS+:MEM_CHANNELS];
				// Trace: src/VX_mem_scheduler.sv:278:13
				assign req_batch_idxs[i * MEM_BATCH_BITS+:MEM_BATCH_BITS] = sv2v_cast_F385D_signed(i);
			end
			// Trace: src/VX_mem_scheduler.sv:280:9
			VX_find_first #(
				.N(MEM_BATCHES),
				.DATAW(MEM_BATCH_BITS),
				.REVERSE(1)
			) find_last(
				.valid_in(req_batch_valids),
				.data_in(req_batch_idxs),
				.data_out(req_batch_idx_last),
				.valid_out()
			);
			// Trace: src/VX_mem_scheduler.sv:290:9
			assign mem_req_valid_s = mem_req_valid_b;
			// Trace: src/VX_mem_scheduler.sv:291:9
			assign req_batch_idx = req_batch_idx_r;
			// Trace: src/VX_mem_scheduler.sv:292:9
			assign req_sent_all = mem_req_ready_b && (req_batch_idx_r == req_batch_idx_last);
			// Trace: src/VX_mem_scheduler.sv:293:9
			assign mem_req_tag_s = {reqq_tag_s, req_batch_idx};
		end
		else begin : g_no_batch
			// Trace: src/VX_mem_scheduler.sv:295:9
			assign mem_req_valid_s = reqq_valid_s;
			// Trace: src/VX_mem_scheduler.sv:296:9
			assign req_batch_idx = 1'sb0;
			// Trace: src/VX_mem_scheduler.sv:297:9
			assign req_sent_all = mem_req_ready_s;
			// Trace: src/VX_mem_scheduler.sv:298:9
			assign mem_req_tag_s = reqq_tag_s;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:300:5
	assign reqq_ready_s = req_sent_all;
	// Trace: src/VX_mem_scheduler.sv:301:5
	wire [(MEM_CHANNELS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] mem_req_flags_u;
	// Trace: src/VX_mem_scheduler.sv:302:5
	VX_elastic_buffer #(
		.DATAW(((MEM_CHANNELS + 1) + (MEM_CHANNELS * (((LINE_SIZE + MEM_ADDR_WIDTH) + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + LINE_WIDTH))) + MEM_TAG_WIDTH),
		.SIZE(((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : 2)),
		.OUT_REG(((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : (MEM_OUT_BUF & 7) - 2))
	) mem_req_buf(
		.clk(clk),
		.reset(reset),
		.valid_in(mem_req_valid_s),
		.ready_in(mem_req_ready_s),
		.data_in({mem_req_mask_s, mem_req_rw_s, mem_req_byteen_s, mem_req_addr_s, mem_req_flags_s, mem_req_data_s, mem_req_tag_s}),
		.data_out({mem_req_mask, mem_req_rw, mem_req_byteen, mem_req_addr, mem_req_flags_u, mem_req_data, mem_req_tag}),
		.valid_out(mem_req_valid),
		.ready_out(mem_req_ready)
	);
	// Trace: src/VX_mem_scheduler.sv:316:5
	generate
		if (FLAGS_WIDTH != 0) begin : g_mem_req_flags
			// Trace: src/VX_mem_scheduler.sv:317:9
			assign mem_req_flags = mem_req_flags_u;
		end
		else begin : g_mem_req_flags_0
			// Trace: src/VX_mem_scheduler.sv:319:9
			assign mem_req_flags = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:321:5
	wire [BATCH_SEL_WIDTH - 1:0] rsp_batch_idx;
	// Trace: src/VX_mem_scheduler.sv:322:5
	generate
		if (CORE_BATCHES > 1) begin : g_rsp_batch_idx
			// Trace: src/VX_mem_scheduler.sv:323:9
			assign rsp_batch_idx = mem_rsp_tag_s[CORE_BATCH_BITS - 1:0];
		end
		else begin : g_rsp_batch_idx_0
			// Trace: src/VX_mem_scheduler.sv:325:9
			assign rsp_batch_idx = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:327:5
	function automatic signed [BATCH_SEL_WIDTH - 1:0] sv2v_cast_397F3_signed;
		input reg signed [BATCH_SEL_WIDTH - 1:0] inp;
		sv2v_cast_397F3_signed = inp;
	endfunction
	generate
		if (CORE_REQS == 1) begin : g_rsp_1
			// Trace: src/VX_mem_scheduler.sv:328:9
			assign crsp_valid = mem_rsp_valid_s;
			// Trace: src/VX_mem_scheduler.sv:329:9
			assign crsp_mask = mem_rsp_mask_s;
			// Trace: src/VX_mem_scheduler.sv:330:9
			assign crsp_sop = 1'b1;
			// Trace: src/VX_mem_scheduler.sv:331:9
			assign crsp_eop = 1'b1;
			// Trace: src/VX_mem_scheduler.sv:332:9
			assign crsp_data = mem_rsp_data_s;
			// Trace: src/VX_mem_scheduler.sv:333:9
			assign mem_rsp_ready_s = crsp_ready;
		end
		else begin : g_rsp_N
			// Trace: src/VX_mem_scheduler.sv:335:9
			reg [(CORE_QUEUE_SIZE * CORE_REQS) - 1:0] rsp_rem_mask;
			// Trace: src/VX_mem_scheduler.sv:336:9
			wire [CORE_REQS - 1:0] rsp_rem_mask_n;
			wire [CORE_REQS - 1:0] curr_mask;
			genvar _gv_r_1;
			for (_gv_r_1 = 0; _gv_r_1 < CORE_REQS; _gv_r_1 = _gv_r_1 + 1) begin : g_curr_mask
				localparam r = _gv_r_1;
				// Trace: src/VX_mem_scheduler.sv:338:13
				localparam i = r / CORE_CHANNELS;
				// Trace: src/VX_mem_scheduler.sv:339:13
				localparam j = r % CORE_CHANNELS;
				// Trace: src/VX_mem_scheduler.sv:340:13
				assign curr_mask[r] = (sv2v_cast_397F3_signed(i) == rsp_batch_idx) && mem_rsp_mask_s[j];
			end
			// Trace: src/VX_mem_scheduler.sv:342:9
			assign rsp_rem_mask_n = rsp_rem_mask[ibuf_raddr * CORE_REQS+:CORE_REQS] & ~curr_mask;
			// Trace: src/VX_mem_scheduler.sv:343:9
			wire mem_rsp_fire_s = mem_rsp_valid_s && mem_rsp_ready_s;
			// Trace: src/VX_mem_scheduler.sv:344:9
			always @(posedge clk) begin
				// Trace: src/VX_mem_scheduler.sv:345:13
				if (ibuf_push)
					// Trace: src/VX_mem_scheduler.sv:346:17
					rsp_rem_mask[ibuf_waddr * CORE_REQS+:CORE_REQS] <= core_req_mask;
				if (mem_rsp_fire_s)
					// Trace: src/VX_mem_scheduler.sv:349:17
					rsp_rem_mask[ibuf_raddr * CORE_REQS+:CORE_REQS] <= rsp_rem_mask_n;
			end
			// Trace: src/VX_mem_scheduler.sv:352:9
			wire rsp_complete = ~(|rsp_rem_mask_n) || (CORE_REQS == 1);
			if (RSP_PARTIAL != 0) begin : g_rsp_partial
				// Trace: src/VX_mem_scheduler.sv:354:13
				reg [CORE_QUEUE_SIZE - 1:0] rsp_sop_r;
				// Trace: src/VX_mem_scheduler.sv:355:13
				always @(posedge clk) begin
					// Trace: src/VX_mem_scheduler.sv:356:17
					if (ibuf_push)
						// Trace: src/VX_mem_scheduler.sv:357:21
						rsp_sop_r[ibuf_waddr] <= 1;
					if (mem_rsp_fire_s)
						// Trace: src/VX_mem_scheduler.sv:360:21
						rsp_sop_r[ibuf_raddr] <= 0;
				end
				// Trace: src/VX_mem_scheduler.sv:363:13
				assign crsp_valid = mem_rsp_valid_s;
				// Trace: src/VX_mem_scheduler.sv:364:13
				assign crsp_mask = curr_mask;
				// Trace: src/VX_mem_scheduler.sv:365:13
				assign crsp_sop = rsp_sop_r[ibuf_raddr];
				genvar _gv_r_2;
				for (_gv_r_2 = 0; _gv_r_2 < CORE_REQS; _gv_r_2 = _gv_r_2 + 1) begin : g_crsp_data
					localparam r = _gv_r_2;
					// Trace: src/VX_mem_scheduler.sv:367:17
					localparam j = r % CORE_CHANNELS;
					// Trace: src/VX_mem_scheduler.sv:368:17
					assign crsp_data[r * WORD_WIDTH+:WORD_WIDTH] = mem_rsp_data_s[j * WORD_WIDTH+:WORD_WIDTH];
				end
				// Trace: src/VX_mem_scheduler.sv:370:13
				assign mem_rsp_ready_s = crsp_ready;
			end
			else begin : g_rsp_full
				// Trace: src/VX_mem_scheduler.sv:372:13
				wire [((CORE_CHANNELS * CORE_BATCHES) * WORD_WIDTH) - 1:0] rsp_store_n;
				// Trace: src/VX_mem_scheduler.sv:373:13
				reg [CORE_REQS - 1:0] rsp_orig_mask [CORE_QUEUE_SIZE - 1:0];
				genvar _gv_i_92;
				for (_gv_i_92 = 0; _gv_i_92 < CORE_CHANNELS; _gv_i_92 = _gv_i_92 + 1) begin : g_rsp_store
					localparam i = _gv_i_92;
					genvar _gv_j_9;
					for (_gv_j_9 = 0; _gv_j_9 < CORE_BATCHES; _gv_j_9 = _gv_j_9 + 1) begin : g_j
						localparam j = _gv_j_9;
						// Trace: src/VX_mem_scheduler.sv:376:21
						reg [WORD_WIDTH - 1:0] rsp_store [0:CORE_QUEUE_SIZE - 1];
						// Trace: src/VX_mem_scheduler.sv:377:21
						wire rsp_wren = (mem_rsp_fire_s && (sv2v_cast_397F3_signed(j) == rsp_batch_idx)) && ((CORE_CHANNELS == 1) || mem_rsp_mask_s[i]);
						// Trace: src/VX_mem_scheduler.sv:380:21
						always @(posedge clk)
							// Trace: src/VX_mem_scheduler.sv:381:25
							if (rsp_wren)
								// Trace: src/VX_mem_scheduler.sv:382:29
								rsp_store[ibuf_raddr] <= mem_rsp_data_s[i * WORD_WIDTH+:WORD_WIDTH];
						// Trace: src/VX_mem_scheduler.sv:385:21
						assign rsp_store_n[((i * CORE_BATCHES) + j) * WORD_WIDTH+:WORD_WIDTH] = (rsp_wren ? mem_rsp_data_s[i * WORD_WIDTH+:WORD_WIDTH] : rsp_store[ibuf_raddr]);
					end
				end
				// Trace: src/VX_mem_scheduler.sv:388:13
				always @(posedge clk)
					// Trace: src/VX_mem_scheduler.sv:389:17
					if (ibuf_push)
						// Trace: src/VX_mem_scheduler.sv:390:21
						rsp_orig_mask[ibuf_waddr] <= core_req_mask;
				// Trace: src/VX_mem_scheduler.sv:393:13
				assign crsp_valid = mem_rsp_valid_s && rsp_complete;
				// Trace: src/VX_mem_scheduler.sv:394:13
				assign crsp_mask = rsp_orig_mask[ibuf_raddr];
				// Trace: src/VX_mem_scheduler.sv:395:13
				assign crsp_sop = 1'b1;
				genvar _gv_r_3;
				for (_gv_r_3 = 0; _gv_r_3 < CORE_REQS; _gv_r_3 = _gv_r_3 + 1) begin : g_crsp_data
					localparam r = _gv_r_3;
					// Trace: src/VX_mem_scheduler.sv:397:17
					localparam i = r / CORE_CHANNELS;
					// Trace: src/VX_mem_scheduler.sv:398:17
					localparam j = r % CORE_CHANNELS;
					// Trace: src/VX_mem_scheduler.sv:399:17
					assign crsp_data[r * WORD_WIDTH+:WORD_WIDTH] = rsp_store_n[((j * CORE_BATCHES) + i) * WORD_WIDTH+:WORD_WIDTH];
				end
				// Trace: src/VX_mem_scheduler.sv:401:13
				assign mem_rsp_ready_s = crsp_ready || ~rsp_complete;
			end
			// Trace: src/VX_mem_scheduler.sv:403:9
			assign crsp_eop = rsp_complete;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:405:5
	generate
		if (UUID_WIDTH != 0) begin : g_crsp_tag
			// Trace: src/VX_mem_scheduler.sv:406:9
			assign crsp_tag = {mem_rsp_tag_s[MEM_TAG_WIDTH - 1-:UUID_WIDTH], ibuf_dout};
		end
		else begin : g_crsp_tag_0
			// Trace: src/VX_mem_scheduler.sv:408:9
			assign crsp_tag = ibuf_dout;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:410:5
	VX_elastic_buffer #(
		.DATAW(((CORE_REQS + 2) + (CORE_REQS * WORD_WIDTH)) + TAG_WIDTH),
		.SIZE(((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : 2)),
		.OUT_REG(((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : (CORE_OUT_BUF & 7) - 2))
	) rsp_buf(
		.clk(clk),
		.reset(reset),
		.valid_in(crsp_valid),
		.ready_in(crsp_ready),
		.data_in({crsp_mask, crsp_sop, crsp_eop, crsp_data, crsp_tag}),
		.data_out({core_rsp_mask, core_rsp_sop, core_rsp_eop, core_rsp_data, core_rsp_tag}),
		.valid_out(core_rsp_valid),
		.ready_out(core_rsp_ready)
	);
endmodule
module VX_pending_size (
	clk,
	reset,
	incr,
	decr,
	empty,
	alm_empty,
	full,
	alm_full,
	size
);
	// Trace: src/VX_pending_size.sv:2:15
	parameter SIZE = 1;
	// Trace: src/VX_pending_size.sv:3:15
	parameter INCRW = 1;
	// Trace: src/VX_pending_size.sv:4:15
	parameter DECRW = 1;
	// Trace: src/VX_pending_size.sv:5:15
	parameter ALM_FULL = SIZE - 1;
	// Trace: src/VX_pending_size.sv:6:15
	parameter ALM_EMPTY = 1;
	// Trace: src/VX_pending_size.sv:7:15
	parameter SIZEW = $clog2(SIZE + 1);
	// Trace: src/VX_pending_size.sv:9:5
	input wire clk;
	// Trace: src/VX_pending_size.sv:10:5
	input wire reset;
	// Trace: src/VX_pending_size.sv:11:5
	input wire [INCRW - 1:0] incr;
	// Trace: src/VX_pending_size.sv:12:5
	input wire [DECRW - 1:0] decr;
	// Trace: src/VX_pending_size.sv:13:5
	output wire empty;
	// Trace: src/VX_pending_size.sv:14:5
	output wire alm_empty;
	// Trace: src/VX_pending_size.sv:15:5
	output wire full;
	// Trace: src/VX_pending_size.sv:16:5
	output wire alm_full;
	// Trace: src/VX_pending_size.sv:17:5
	output wire [SIZEW - 1:0] size;
	// Trace: src/VX_pending_size.sv:19:5
	function automatic signed [SIZEW - 1:0] sv2v_cast_33A93_signed;
		input reg signed [SIZEW - 1:0] inp;
		sv2v_cast_33A93_signed = inp;
	endfunction
	generate
		if (SIZE == 1) begin : g_size_eq1
			// Trace: src/VX_pending_size.sv:20:9
			reg size_r;
			// Trace: src/VX_pending_size.sv:21:9
			always @(posedge clk)
				// Trace: src/VX_pending_size.sv:22:13
				if (reset)
					// Trace: src/VX_pending_size.sv:23:17
					size_r <= 1'sb0;
				else
					// Trace: src/VX_pending_size.sv:25:17
					if (incr) begin
						begin
							// Trace: src/VX_pending_size.sv:26:21
							if (~decr)
								// Trace: src/VX_pending_size.sv:27:25
								size_r <= 1;
						end
					end
					else if (decr)
						// Trace: src/VX_pending_size.sv:30:21
						size_r <= 1'sb0;
			// Trace: src/VX_pending_size.sv:34:9
			assign empty = size_r == 0;
			// Trace: src/VX_pending_size.sv:35:9
			assign full = size_r != 0;
			// Trace: src/VX_pending_size.sv:36:9
			assign alm_empty = 1'b1;
			// Trace: src/VX_pending_size.sv:37:9
			assign alm_full = 1'b1;
			// Trace: src/VX_pending_size.sv:38:9
			assign size = size_r;
		end
		else begin : g_size_gt1
			// Trace: src/VX_pending_size.sv:40:9
			reg empty_r;
			reg alm_empty_r;
			// Trace: src/VX_pending_size.sv:41:9
			reg full_r;
			reg alm_full_r;
			if ((INCRW != 1) || (DECRW != 1)) begin : g_wide_step
				// Trace: src/VX_pending_size.sv:43:13
				localparam DELTAW = (SIZEW < ((INCRW > DECRW ? INCRW : DECRW) + 1) ? SIZEW : (INCRW > DECRW ? INCRW : DECRW) + 1);
				// Trace: src/VX_pending_size.sv:44:13
				wire [SIZEW - 1:0] size_n;
				reg [SIZEW - 1:0] size_r;
				// Trace: src/VX_pending_size.sv:45:13
				function automatic [DELTAW - 1:0] sv2v_cast_B4011;
					input reg [DELTAW - 1:0] inp;
					sv2v_cast_B4011 = inp;
				endfunction
				wire [DELTAW - 1:0] delta = sv2v_cast_B4011(incr) - sv2v_cast_B4011(decr);
				// Trace: src/VX_pending_size.sv:46:13
				assign size_n = $signed(size_r) + sv2v_cast_33A93_signed($signed(delta));
				// Trace: src/VX_pending_size.sv:47:13
				always @(posedge clk)
					// Trace: src/VX_pending_size.sv:48:17
					if (reset) begin
						// Trace: src/VX_pending_size.sv:49:21
						empty_r <= 1;
						// Trace: src/VX_pending_size.sv:50:21
						full_r <= 0;
						// Trace: src/VX_pending_size.sv:51:21
						alm_empty_r <= 1;
						// Trace: src/VX_pending_size.sv:52:21
						alm_full_r <= 0;
						// Trace: src/VX_pending_size.sv:53:21
						size_r <= 1'sb0;
					end
					else begin
						// Trace: src/VX_pending_size.sv:55:21
						// Trace: src/VX_pending_size.sv:57:21
						empty_r <= size_n == sv2v_cast_33A93_signed(0);
						// Trace: src/VX_pending_size.sv:58:21
						full_r <= size_n == sv2v_cast_33A93_signed(SIZE);
						// Trace: src/VX_pending_size.sv:59:21
						alm_empty_r <= size_n <= sv2v_cast_33A93_signed(ALM_EMPTY);
						// Trace: src/VX_pending_size.sv:60:21
						alm_full_r <= size_n >= sv2v_cast_33A93_signed(ALM_FULL);
						// Trace: src/VX_pending_size.sv:61:21
						size_r <= size_n;
					end
				// Trace: src/VX_pending_size.sv:64:13
				assign size = size_r;
			end
			else begin : g_single_step
				// Trace: src/VX_pending_size.sv:66:13
				localparam ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
				// Trace: src/VX_pending_size.sv:67:13
				reg [ADDRW - 1:0] used_r;
				// Trace: src/VX_pending_size.sv:68:13
				function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
					input reg signed [ADDRW - 1:0] inp;
					sv2v_cast_8BB5D_signed = inp;
				endfunction
				wire is_alm_empty = used_r == sv2v_cast_8BB5D_signed(ALM_EMPTY);
				// Trace: src/VX_pending_size.sv:69:13
				wire is_alm_empty_n = used_r == sv2v_cast_8BB5D_signed(ALM_EMPTY + 1);
				// Trace: src/VX_pending_size.sv:70:13
				wire is_alm_full = used_r == sv2v_cast_8BB5D_signed(ALM_FULL);
				// Trace: src/VX_pending_size.sv:71:13
				wire is_alm_full_n = used_r == sv2v_cast_8BB5D_signed(ALM_FULL - 1);
				// Trace: src/VX_pending_size.sv:72:13
				always @(posedge clk)
					// Trace: src/VX_pending_size.sv:73:17
					if (reset) begin
						// Trace: src/VX_pending_size.sv:74:21
						alm_empty_r <= 1;
						// Trace: src/VX_pending_size.sv:75:21
						alm_full_r <= 0;
					end
					else
						// Trace: src/VX_pending_size.sv:77:21
						if (incr) begin
							begin
								// Trace: src/VX_pending_size.sv:78:25
								if (~decr) begin
									// Trace: src/VX_pending_size.sv:79:29
									if (is_alm_empty)
										// Trace: src/VX_pending_size.sv:80:33
										alm_empty_r <= 0;
									if (is_alm_full_n)
										// Trace: src/VX_pending_size.sv:82:33
										alm_full_r <= 1;
								end
							end
						end
						else if (decr) begin
							// Trace: src/VX_pending_size.sv:85:25
							if (is_alm_full)
								// Trace: src/VX_pending_size.sv:86:29
								alm_full_r <= 0;
							if (is_alm_empty_n)
								// Trace: src/VX_pending_size.sv:88:29
								alm_empty_r <= 1;
						end
				if (SIZE > 2) begin : g_size_gt2
					// Trace: src/VX_pending_size.sv:93:17
					function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
						input reg signed [ADDRW - 1:0] inp;
						sv2v_cast_8BB5D_signed = inp;
					endfunction
					wire is_empty_n = used_r == sv2v_cast_8BB5D_signed(1);
					// Trace: src/VX_pending_size.sv:94:17
					wire is_full_n = used_r == sv2v_cast_8BB5D_signed(SIZE - 1);
					// Trace: src/VX_pending_size.sv:95:17
					wire [1:0] delta = {~incr & decr, incr ^ decr};
					// Trace: src/VX_pending_size.sv:96:17
					always @(posedge clk)
						// Trace: src/VX_pending_size.sv:97:21
						if (reset) begin
							// Trace: src/VX_pending_size.sv:98:25
							empty_r <= 1;
							// Trace: src/VX_pending_size.sv:99:25
							full_r <= 0;
							// Trace: src/VX_pending_size.sv:100:25
							used_r <= 1'sb0;
						end
						else begin
							// Trace: src/VX_pending_size.sv:102:25
							if (incr) begin
								begin
									// Trace: src/VX_pending_size.sv:103:29
									if (~decr) begin
										// Trace: src/VX_pending_size.sv:104:33
										empty_r <= 0;
										// Trace: src/VX_pending_size.sv:105:33
										if (is_full_n)
											// Trace: src/VX_pending_size.sv:106:37
											full_r <= 1;
									end
								end
							end
							else if (decr) begin
								// Trace: src/VX_pending_size.sv:109:29
								full_r <= 0;
								// Trace: src/VX_pending_size.sv:110:29
								if (is_empty_n)
									// Trace: src/VX_pending_size.sv:111:33
									empty_r <= 1;
							end
							// Trace: src/VX_pending_size.sv:113:25
							begin : sv2v_autoblock_1
								reg signed [ADDRW - 1:0] sv2v_tmp_cast;
								sv2v_tmp_cast = $signed(delta);
								used_r <= $signed(used_r) + sv2v_tmp_cast;
							end
						end
				end
				else begin : g_size_eq2
					// Trace: src/VX_pending_size.sv:117:17
					always @(posedge clk)
						// Trace: src/VX_pending_size.sv:118:21
						if (reset) begin
							// Trace: src/VX_pending_size.sv:119:25
							empty_r <= 1;
							// Trace: src/VX_pending_size.sv:120:25
							full_r <= 0;
							// Trace: src/VX_pending_size.sv:121:25
							used_r <= 1'sb0;
						end
						else begin
							// Trace: src/VX_pending_size.sv:123:25
							empty_r <= (empty_r & ~incr) | ((~full_r & decr) & ~incr);
							// Trace: src/VX_pending_size.sv:124:25
							full_r <= ((~empty_r & incr) & ~decr) | (full_r & ~(decr ^ incr));
							// Trace: src/VX_pending_size.sv:125:25
							used_r <= used_r ^ (incr ^ decr);
						end
				end
				if (SIZE > 1) begin : g_sizeN
					if (SIZEW > ADDRW) begin : g_not_log2
						// Trace: src/VX_pending_size.sv:131:21
						assign size = {full_r, used_r};
					end
					else begin : g_log2
						// Trace: src/VX_pending_size.sv:133:21
						assign size = used_r;
					end
				end
				else begin : g_size1
					// Trace: src/VX_pending_size.sv:136:17
					assign size = full_r;
				end
			end
			// Trace: src/VX_pending_size.sv:139:9
			assign empty = empty_r;
			// Trace: src/VX_pending_size.sv:140:9
			assign full = full_r;
			// Trace: src/VX_pending_size.sv:141:9
			assign alm_empty = alm_empty_r;
			// Trace: src/VX_pending_size.sv:142:9
			assign alm_full = alm_full_r;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_ibuffer
// removed module with interface ports: VX_lsu_unit
// removed module with interface ports: VX_lmem_switch
// removed module with interface ports: VX_dispatch_unit
// removed interface: VX_fpu_csr_if
// removed interface: VX_ibuffer_if
module VX_matrix_arbiter (
	clk,
	reset,
	requests,
	grant_index,
	grant_onehot,
	grant_valid,
	grant_ready
);
	// Trace: src/VX_matrix_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_matrix_arbiter.sv:3:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_matrix_arbiter.sv:5:5
	input wire clk;
	// Trace: src/VX_matrix_arbiter.sv:6:5
	input wire reset;
	// Trace: src/VX_matrix_arbiter.sv:7:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_matrix_arbiter.sv:8:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_matrix_arbiter.sv:9:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_matrix_arbiter.sv:10:5
	output wire grant_valid;
	// Trace: src/VX_matrix_arbiter.sv:11:5
	input wire grant_ready;
	// Trace: src/VX_matrix_arbiter.sv:13:5
	generate
		if (NUM_REQS == 1) begin : g_passthru
			// Trace: src/VX_matrix_arbiter.sv:14:9
			assign grant_index = 1'sb0;
			// Trace: src/VX_matrix_arbiter.sv:15:9
			assign grant_onehot = requests;
			// Trace: src/VX_matrix_arbiter.sv:16:9
			assign grant_valid = requests[0];
		end
		else begin : g_arbiter
			// Trace: src/VX_matrix_arbiter.sv:18:9
			reg [NUM_REQS - 1:1] state [NUM_REQS - 1:0];
			// Trace: src/VX_matrix_arbiter.sv:19:9
			wire [NUM_REQS - 1:0] pri [NUM_REQS - 1:0];
			// Trace: src/VX_matrix_arbiter.sv:20:9
			wire [NUM_REQS - 1:0] grant;
			genvar _gv_r_4;
			for (_gv_r_4 = 0; _gv_r_4 < NUM_REQS; _gv_r_4 = _gv_r_4 + 1) begin : g_pri_r
				localparam r = _gv_r_4;
				genvar _gv_c_1;
				for (_gv_c_1 = 0; _gv_c_1 < NUM_REQS; _gv_c_1 = _gv_c_1 + 1) begin : g_pri_c
					localparam c = _gv_c_1;
					if (r > c) begin : g_row
						// Trace: src/VX_matrix_arbiter.sv:24:21
						assign pri[r][c] = requests[c] && state[c][r];
					end
					else if (r < c) begin : g_col
						// Trace: src/VX_matrix_arbiter.sv:26:21
						assign pri[r][c] = requests[c] && !state[r][c];
					end
					else begin : g_equal
						// Trace: src/VX_matrix_arbiter.sv:28:21
						assign pri[r][c] = 0;
					end
				end
			end
			genvar _gv_r_5;
			for (_gv_r_5 = 0; _gv_r_5 < NUM_REQS; _gv_r_5 = _gv_r_5 + 1) begin : g_grant
				localparam r = _gv_r_5;
				// Trace: src/VX_matrix_arbiter.sv:33:13
				assign grant[r] = requests[r] && ~(|pri[r]);
			end
			genvar _gv_r_6;
			for (_gv_r_6 = 0; _gv_r_6 < NUM_REQS; _gv_r_6 = _gv_r_6 + 1) begin : g_state_r
				localparam r = _gv_r_6;
				genvar _gv_c_2;
				for (_gv_c_2 = r + 1; _gv_c_2 < NUM_REQS; _gv_c_2 = _gv_c_2 + 1) begin : g_state_c
					localparam c = _gv_c_2;
					// Trace: src/VX_matrix_arbiter.sv:37:17
					always @(posedge clk)
						// Trace: src/VX_matrix_arbiter.sv:38:21
						if (reset)
							// Trace: src/VX_matrix_arbiter.sv:39:25
							state[r][c] <= 1'sb0;
						else if (grant_ready)
							// Trace: src/VX_matrix_arbiter.sv:41:25
							state[r][c] <= (state[r][c] || grant[c]) && ~grant[r];
				end
			end
			// Trace: src/VX_matrix_arbiter.sv:46:9
			assign grant_onehot = grant;
			// Trace: src/VX_matrix_arbiter.sv:47:9
			VX_onehot_encoder #(.N(NUM_REQS)) encoder(
				.data_in(grant_onehot),
				.data_out(grant_index),
				.valid_out(grant_valid)
			);
		end
	endgenerate
endmodule
module VX_mem_coalescer (
	clk,
	reset,
	in_req_valid,
	in_req_rw,
	in_req_mask,
	in_req_byteen,
	in_req_addr,
	in_req_flags,
	in_req_data,
	in_req_tag,
	in_req_ready,
	in_rsp_valid,
	in_rsp_mask,
	in_rsp_data,
	in_rsp_tag,
	in_rsp_ready,
	out_req_valid,
	out_req_rw,
	out_req_mask,
	out_req_byteen,
	out_req_addr,
	out_req_flags,
	out_req_data,
	out_req_tag,
	out_req_ready,
	out_rsp_valid,
	out_rsp_mask,
	out_rsp_data,
	out_rsp_tag,
	out_rsp_ready
);
	// Trace: src/VX_mem_coalescer.sv:2:15
	parameter INSTANCE_ID = "";
	// Trace: src/VX_mem_coalescer.sv:3:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_mem_coalescer.sv:4:15
	parameter ADDR_WIDTH = 32;
	// Trace: src/VX_mem_coalescer.sv:5:15
	parameter FLAGS_WIDTH = 0;
	// Trace: src/VX_mem_coalescer.sv:6:15
	parameter DATA_IN_SIZE = 4;
	// Trace: src/VX_mem_coalescer.sv:7:15
	parameter DATA_OUT_SIZE = 64;
	// Trace: src/VX_mem_coalescer.sv:8:15
	parameter TAG_WIDTH = 8;
	// Trace: src/VX_mem_coalescer.sv:9:15
	parameter UUID_WIDTH = 0;
	// Trace: src/VX_mem_coalescer.sv:10:15
	parameter QUEUE_SIZE = 8;
	// Trace: src/VX_mem_coalescer.sv:11:15
	parameter DATA_IN_WIDTH = DATA_IN_SIZE * 8;
	// Trace: src/VX_mem_coalescer.sv:12:15
	parameter DATA_OUT_WIDTH = DATA_OUT_SIZE * 8;
	// Trace: src/VX_mem_coalescer.sv:13:15
	parameter DATA_RATIO = DATA_OUT_SIZE / DATA_IN_SIZE;
	// Trace: src/VX_mem_coalescer.sv:14:15
	parameter DATA_RATIO_W = (DATA_RATIO > 1 ? $clog2(DATA_RATIO) : 1);
	// Trace: src/VX_mem_coalescer.sv:15:15
	parameter OUT_REQS = NUM_REQS / DATA_RATIO;
	// Trace: src/VX_mem_coalescer.sv:16:15
	parameter OUT_ADDR_WIDTH = ADDR_WIDTH - DATA_RATIO_W;
	// Trace: src/VX_mem_coalescer.sv:17:15
	parameter QUEUE_ADDRW = $clog2(QUEUE_SIZE);
	// Trace: src/VX_mem_coalescer.sv:18:15
	parameter OUT_TAG_WIDTH = UUID_WIDTH + QUEUE_ADDRW;
	// Trace: src/VX_mem_coalescer.sv:20:5
	input wire clk;
	// Trace: src/VX_mem_coalescer.sv:21:5
	input wire reset;
	// Trace: src/VX_mem_coalescer.sv:22:5
	input wire in_req_valid;
	// Trace: src/VX_mem_coalescer.sv:23:5
	input wire in_req_rw;
	// Trace: src/VX_mem_coalescer.sv:24:5
	input wire [NUM_REQS - 1:0] in_req_mask;
	// Trace: src/VX_mem_coalescer.sv:25:5
	input wire [(NUM_REQS * DATA_IN_SIZE) - 1:0] in_req_byteen;
	// Trace: src/VX_mem_coalescer.sv:26:5
	input wire [(NUM_REQS * ADDR_WIDTH) - 1:0] in_req_addr;
	// Trace: src/VX_mem_coalescer.sv:27:5
	input wire [(NUM_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] in_req_flags;
	// Trace: src/VX_mem_coalescer.sv:28:5
	input wire [(NUM_REQS * DATA_IN_WIDTH) - 1:0] in_req_data;
	// Trace: src/VX_mem_coalescer.sv:29:5
	input wire [TAG_WIDTH - 1:0] in_req_tag;
	// Trace: src/VX_mem_coalescer.sv:30:5
	output wire in_req_ready;
	// Trace: src/VX_mem_coalescer.sv:31:5
	output wire in_rsp_valid;
	// Trace: src/VX_mem_coalescer.sv:32:5
	output wire [NUM_REQS - 1:0] in_rsp_mask;
	// Trace: src/VX_mem_coalescer.sv:33:5
	output wire [(NUM_REQS * DATA_IN_WIDTH) - 1:0] in_rsp_data;
	// Trace: src/VX_mem_coalescer.sv:34:5
	output wire [TAG_WIDTH - 1:0] in_rsp_tag;
	// Trace: src/VX_mem_coalescer.sv:35:5
	input wire in_rsp_ready;
	// Trace: src/VX_mem_coalescer.sv:36:5
	output wire out_req_valid;
	// Trace: src/VX_mem_coalescer.sv:37:5
	output wire out_req_rw;
	// Trace: src/VX_mem_coalescer.sv:38:5
	output wire [OUT_REQS - 1:0] out_req_mask;
	// Trace: src/VX_mem_coalescer.sv:39:5
	output wire [(OUT_REQS * DATA_OUT_SIZE) - 1:0] out_req_byteen;
	// Trace: src/VX_mem_coalescer.sv:40:5
	output wire [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] out_req_addr;
	// Trace: src/VX_mem_coalescer.sv:41:5
	output wire [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] out_req_flags;
	// Trace: src/VX_mem_coalescer.sv:42:5
	output wire [(OUT_REQS * DATA_OUT_WIDTH) - 1:0] out_req_data;
	// Trace: src/VX_mem_coalescer.sv:43:5
	output wire [OUT_TAG_WIDTH - 1:0] out_req_tag;
	// Trace: src/VX_mem_coalescer.sv:44:5
	input wire out_req_ready;
	// Trace: src/VX_mem_coalescer.sv:45:5
	input wire out_rsp_valid;
	// Trace: src/VX_mem_coalescer.sv:46:5
	input wire [OUT_REQS - 1:0] out_rsp_mask;
	// Trace: src/VX_mem_coalescer.sv:47:5
	input wire [(OUT_REQS * DATA_OUT_WIDTH) - 1:0] out_rsp_data;
	// Trace: src/VX_mem_coalescer.sv:48:5
	input wire [OUT_TAG_WIDTH - 1:0] out_rsp_tag;
	// Trace: src/VX_mem_coalescer.sv:49:5
	output wire out_rsp_ready;
	// Trace: src/VX_mem_coalescer.sv:51:5
	localparam TAG_ID_WIDTH = TAG_WIDTH - UUID_WIDTH;
	// Trace: src/VX_mem_coalescer.sv:52:5
	localparam IBUF_DATA_WIDTH = (TAG_ID_WIDTH + NUM_REQS) + (NUM_REQS * DATA_RATIO_W);
	// Trace: src/VX_mem_coalescer.sv:53:5
	localparam STATE_WAIT = 0;
	// Trace: src/VX_mem_coalescer.sv:54:5
	localparam STATE_SEND = 1;
	// Trace: src/VX_mem_coalescer.sv:55:5
	wire state_r;
	reg state_n;
	// Trace: src/VX_mem_coalescer.sv:56:5
	wire out_req_valid_r;
	reg out_req_valid_n;
	// Trace: src/VX_mem_coalescer.sv:57:5
	wire out_req_rw_r;
	reg out_req_rw_n;
	// Trace: src/VX_mem_coalescer.sv:58:5
	wire [OUT_REQS - 1:0] out_req_mask_r;
	reg [OUT_REQS - 1:0] out_req_mask_n;
	// Trace: src/VX_mem_coalescer.sv:59:5
	wire [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] out_req_addr_r;
	reg [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] out_req_addr_n;
	// Trace: src/VX_mem_coalescer.sv:60:5
	wire [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] out_req_flags_r;
	reg [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] out_req_flags_n;
	// Trace: src/VX_mem_coalescer.sv:61:5
	wire [((OUT_REQS * DATA_RATIO) * DATA_IN_SIZE) - 1:0] out_req_byteen_r;
	reg [((OUT_REQS * DATA_RATIO) * DATA_IN_SIZE) - 1:0] out_req_byteen_n;
	// Trace: src/VX_mem_coalescer.sv:62:5
	wire [((OUT_REQS * DATA_RATIO) * DATA_IN_WIDTH) - 1:0] out_req_data_r;
	reg [((OUT_REQS * DATA_RATIO) * DATA_IN_WIDTH) - 1:0] out_req_data_n;
	// Trace: src/VX_mem_coalescer.sv:63:5
	wire [OUT_TAG_WIDTH - 1:0] out_req_tag_r;
	reg [OUT_TAG_WIDTH - 1:0] out_req_tag_n;
	// Trace: src/VX_mem_coalescer.sv:64:5
	reg in_req_ready_n;
	// Trace: src/VX_mem_coalescer.sv:65:5
	wire ibuf_push;
	// Trace: src/VX_mem_coalescer.sv:66:5
	wire ibuf_pop;
	// Trace: src/VX_mem_coalescer.sv:67:5
	wire [QUEUE_ADDRW - 1:0] ibuf_waddr;
	// Trace: src/VX_mem_coalescer.sv:68:5
	wire [QUEUE_ADDRW - 1:0] ibuf_raddr;
	// Trace: src/VX_mem_coalescer.sv:69:5
	wire ibuf_full;
	// Trace: src/VX_mem_coalescer.sv:70:5
	wire ibuf_empty;
	// Trace: src/VX_mem_coalescer.sv:71:5
	wire [IBUF_DATA_WIDTH - 1:0] ibuf_din;
	// Trace: src/VX_mem_coalescer.sv:72:5
	wire [IBUF_DATA_WIDTH - 1:0] ibuf_dout;
	// Trace: src/VX_mem_coalescer.sv:73:5
	wire [OUT_REQS - 1:0] batch_valid_r;
	wire [OUT_REQS - 1:0] batch_valid_n;
	// Trace: src/VX_mem_coalescer.sv:74:5
	wire [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] seed_addr_r;
	wire [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] seed_addr_n;
	// Trace: src/VX_mem_coalescer.sv:75:5
	wire [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] seed_flags_r;
	wire [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] seed_flags_n;
	// Trace: src/VX_mem_coalescer.sv:76:5
	wire [NUM_REQS - 1:0] addr_matches_r;
	wire [NUM_REQS - 1:0] addr_matches_n;
	// Trace: src/VX_mem_coalescer.sv:77:5
	wire [NUM_REQS - 1:0] req_rem_mask_r;
	reg [NUM_REQS - 1:0] req_rem_mask_n;
	// Trace: src/VX_mem_coalescer.sv:78:5
	wire [(NUM_REQS * DATA_RATIO_W) - 1:0] in_addr_offset;
	// Trace: src/VX_mem_coalescer.sv:79:5
	genvar _gv_i_101;
	generate
		for (_gv_i_101 = 0; _gv_i_101 < NUM_REQS; _gv_i_101 = _gv_i_101 + 1) begin : g_in_addr_offset
			localparam i = _gv_i_101;
			// Trace: src/VX_mem_coalescer.sv:80:9
			assign in_addr_offset[i * DATA_RATIO_W+:DATA_RATIO_W] = in_req_addr[(i * ADDR_WIDTH) + (DATA_RATIO_W - 1)-:DATA_RATIO_W];
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:82:5
	genvar _gv_i_102;
	generate
		for (_gv_i_102 = 0; _gv_i_102 < OUT_REQS; _gv_i_102 = _gv_i_102 + 1) begin : g_seed_gen
			localparam i = _gv_i_102;
			// Trace: src/VX_mem_coalescer.sv:83:9
			wire [DATA_RATIO - 1:0] batch_mask;
			// Trace: src/VX_mem_coalescer.sv:84:9
			wire [DATA_RATIO_W - 1:0] batch_idx;
			// Trace: src/VX_mem_coalescer.sv:85:9
			assign batch_mask = in_req_mask[i * DATA_RATIO+:DATA_RATIO] & req_rem_mask_r[i * DATA_RATIO+:DATA_RATIO];
			// Trace: src/VX_mem_coalescer.sv:86:9
			VX_priority_encoder #(.N(DATA_RATIO)) priority_encoder(
				.data_in(batch_mask),
				.index_out(batch_idx),
				.onehot_out(),
				.valid_out(batch_valid_n[i])
			);
			// Trace: src/VX_mem_coalescer.sv:94:9
			wire [(DATA_RATIO * OUT_ADDR_WIDTH) - 1:0] addr_base;
			genvar _gv_j_11;
			for (_gv_j_11 = 0; _gv_j_11 < DATA_RATIO; _gv_j_11 = _gv_j_11 + 1) begin : g_addr_base
				localparam j = _gv_j_11;
				// Trace: src/VX_mem_coalescer.sv:96:13
				assign addr_base[j * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH] = in_req_addr[(((DATA_RATIO * i) + j) * ADDR_WIDTH) + ((ADDR_WIDTH - 1) >= DATA_RATIO_W ? ADDR_WIDTH - 1 : ((ADDR_WIDTH - 1) + ((ADDR_WIDTH - 1) >= DATA_RATIO_W ? ((ADDR_WIDTH - 1) - DATA_RATIO_W) + 1 : (DATA_RATIO_W - (ADDR_WIDTH - 1)) + 1)) - 1)-:((ADDR_WIDTH - 1) >= DATA_RATIO_W ? ((ADDR_WIDTH - 1) - DATA_RATIO_W) + 1 : (DATA_RATIO_W - (ADDR_WIDTH - 1)) + 1)];
			end
			// Trace: src/VX_mem_coalescer.sv:98:9
			wire [(DATA_RATIO * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] req_flags;
			genvar _gv_j_12;
			for (_gv_j_12 = 0; _gv_j_12 < DATA_RATIO; _gv_j_12 = _gv_j_12 + 1) begin : g_req_flags
				localparam j = _gv_j_12;
				// Trace: src/VX_mem_coalescer.sv:100:13
				assign req_flags[j * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)] = in_req_flags[((DATA_RATIO * i) + j) * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)];
			end
			// Trace: src/VX_mem_coalescer.sv:102:9
			assign seed_addr_n[i * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH] = addr_base[batch_idx * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH];
			// Trace: src/VX_mem_coalescer.sv:103:9
			assign seed_flags_n[i * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)] = req_flags[batch_idx * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)];
			genvar _gv_j_13;
			for (_gv_j_13 = 0; _gv_j_13 < DATA_RATIO; _gv_j_13 = _gv_j_13 + 1) begin : g_addr_matches_n
				localparam j = _gv_j_13;
				// Trace: src/VX_mem_coalescer.sv:105:13
				assign addr_matches_n[(i * DATA_RATIO) + j] = addr_base[j * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH] == seed_addr_n[i * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH];
			end
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:108:5
	wire [NUM_REQS - 1:0] current_pmask = in_req_mask & addr_matches_r;
	// Trace: src/VX_mem_coalescer.sv:109:5
	wire [((OUT_REQS * DATA_RATIO) * DATA_IN_SIZE) - 1:0] req_byteen_merged;
	// Trace: src/VX_mem_coalescer.sv:110:5
	wire [((OUT_REQS * DATA_RATIO) * DATA_IN_WIDTH) - 1:0] req_data_merged;
	// Trace: src/VX_mem_coalescer.sv:111:5
	genvar _gv_i_103;
	generate
		for (_gv_i_103 = 0; _gv_i_103 < OUT_REQS; _gv_i_103 = _gv_i_103 + 1) begin : g_data_merged
			localparam i = _gv_i_103;
			// Trace: src/VX_mem_coalescer.sv:112:9
			reg [(DATA_RATIO * DATA_IN_SIZE) - 1:0] byteen_merged;
			// Trace: src/VX_mem_coalescer.sv:113:9
			reg [(DATA_RATIO * DATA_IN_WIDTH) - 1:0] data_merged;
			// Trace: src/VX_mem_coalescer.sv:114:9
			always @(*) begin
				// Trace: src/VX_mem_coalescer.sv:115:13
				byteen_merged = 1'sb0;
				// Trace: src/VX_mem_coalescer.sv:116:13
				data_merged = 1'sbx;
				// Trace: src/VX_mem_coalescer.sv:117:13
				begin : sv2v_autoblock_1
					// Trace: src/VX_mem_coalescer.sv:117:18
					integer j;
					// Trace: src/VX_mem_coalescer.sv:117:18
					for (j = 0; j < DATA_RATIO; j = j + 1)
						begin
							// Trace: src/VX_mem_coalescer.sv:118:17
							begin : sv2v_autoblock_2
								// Trace: src/VX_mem_coalescer.sv:118:22
								integer k;
								// Trace: src/VX_mem_coalescer.sv:118:22
								for (k = 0; k < DATA_IN_SIZE; k = k + 1)
									begin
										// Trace: src/VX_mem_coalescer.sv:119:21
										if (current_pmask[(i * DATA_RATIO) + j] && in_req_byteen[(((DATA_RATIO * i) + j) * DATA_IN_SIZE) + k]) begin
											// Trace: src/VX_mem_coalescer.sv:120:25
											byteen_merged[(in_addr_offset[((DATA_RATIO * i) + j) * DATA_RATIO_W+:DATA_RATIO_W] * DATA_IN_SIZE) + k] = 1'b1;
											// Trace: src/VX_mem_coalescer.sv:121:25
											data_merged[(in_addr_offset[((DATA_RATIO * i) + j) * DATA_RATIO_W+:DATA_RATIO_W] * DATA_IN_WIDTH) + (k * 8)+:8] = in_req_data[(((DATA_RATIO * i) + j) * DATA_IN_WIDTH) + (k * 8)+:8];
										end
									end
							end
						end
				end
			end
			// Trace: src/VX_mem_coalescer.sv:126:9
			assign req_byteen_merged[DATA_IN_SIZE * (i * DATA_RATIO)+:DATA_IN_SIZE * DATA_RATIO] = byteen_merged;
			// Trace: src/VX_mem_coalescer.sv:127:9
			assign req_data_merged[DATA_IN_WIDTH * (i * DATA_RATIO)+:DATA_IN_WIDTH * DATA_RATIO] = data_merged;
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:129:5
	wire is_last_batch = ~(|((in_req_mask & ~addr_matches_r) & req_rem_mask_r));
	// Trace: src/VX_mem_coalescer.sv:130:5
	wire out_req_fire = out_req_valid && out_req_ready;
	// Trace: src/VX_mem_coalescer.sv:131:5
	always @(*) begin
		// Trace: src/VX_mem_coalescer.sv:132:9
		state_n = state_r;
		// Trace: src/VX_mem_coalescer.sv:133:9
		out_req_valid_n = out_req_valid_r;
		// Trace: src/VX_mem_coalescer.sv:134:9
		out_req_mask_n = out_req_mask_r;
		// Trace: src/VX_mem_coalescer.sv:135:9
		out_req_rw_n = out_req_rw_r;
		// Trace: src/VX_mem_coalescer.sv:136:9
		out_req_addr_n = out_req_addr_r;
		// Trace: src/VX_mem_coalescer.sv:137:9
		out_req_flags_n = out_req_flags_r;
		// Trace: src/VX_mem_coalescer.sv:138:9
		out_req_byteen_n = out_req_byteen_r;
		// Trace: src/VX_mem_coalescer.sv:139:9
		out_req_data_n = out_req_data_r;
		// Trace: src/VX_mem_coalescer.sv:140:9
		out_req_tag_n = out_req_tag_r;
		// Trace: src/VX_mem_coalescer.sv:141:9
		req_rem_mask_n = req_rem_mask_r;
		// Trace: src/VX_mem_coalescer.sv:142:9
		in_req_ready_n = 0;
		// Trace: src/VX_mem_coalescer.sv:143:9
		case (state_r)
			STATE_WAIT: begin
				// Trace: src/VX_mem_coalescer.sv:145:13
				if (out_req_fire)
					// Trace: src/VX_mem_coalescer.sv:146:17
					out_req_valid_n = 0;
				if ((in_req_valid && ~out_req_valid_n) && ~ibuf_full)
					// Trace: src/VX_mem_coalescer.sv:149:17
					state_n = STATE_SEND;
			end
			default: begin
				// Trace: src/VX_mem_coalescer.sv:153:13
				state_n = STATE_WAIT;
				// Trace: src/VX_mem_coalescer.sv:154:13
				out_req_valid_n = 1;
				// Trace: src/VX_mem_coalescer.sv:155:13
				out_req_mask_n = batch_valid_r;
				// Trace: src/VX_mem_coalescer.sv:156:13
				out_req_rw_n = in_req_rw;
				// Trace: src/VX_mem_coalescer.sv:157:13
				out_req_addr_n = seed_addr_r;
				// Trace: src/VX_mem_coalescer.sv:158:13
				out_req_flags_n = seed_flags_r;
				// Trace: src/VX_mem_coalescer.sv:159:13
				out_req_byteen_n = req_byteen_merged;
				// Trace: src/VX_mem_coalescer.sv:160:13
				out_req_data_n = req_data_merged;
				// Trace: src/VX_mem_coalescer.sv:161:13
				out_req_tag_n = {in_req_tag[TAG_WIDTH - 1-:UUID_WIDTH], ibuf_waddr};
				// Trace: src/VX_mem_coalescer.sv:162:13
				req_rem_mask_n = (is_last_batch ? {NUM_REQS {1'sb1}} : req_rem_mask_r & ~current_pmask);
				// Trace: src/VX_mem_coalescer.sv:163:13
				in_req_ready_n = is_last_batch;
			end
		endcase
	end
	// Trace: src/VX_mem_coalescer.sv:167:5
	VX_pipe_register #(
		.DATAW(((((1 + NUM_REQS) + 2) + NUM_REQS) + (OUT_REQS * ((((((2 + OUT_ADDR_WIDTH) + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + OUT_ADDR_WIDTH) + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + DATA_OUT_SIZE) + DATA_OUT_WIDTH))) + OUT_TAG_WIDTH),
		.RESETW((1 + NUM_REQS) + 1),
		.INIT_VALUE({1'b0, {NUM_REQS {1'b1}}, 1'b0})
	) pipe_reg(
		.clk(clk),
		.reset(reset),
		.enable(1'b1),
		.data_in({state_n, req_rem_mask_n, out_req_valid_n, out_req_rw_n, addr_matches_n, batch_valid_n, out_req_mask_n, seed_addr_n, seed_flags_n, out_req_addr_n, out_req_flags_n, out_req_byteen_n, out_req_data_n, out_req_tag_n}),
		.data_out({state_r, req_rem_mask_r, out_req_valid_r, out_req_rw_r, addr_matches_r, batch_valid_r, out_req_mask_r, seed_addr_r, seed_flags_r, out_req_addr_r, out_req_flags_r, out_req_byteen_r, out_req_data_r, out_req_tag_r})
	);
	// Trace: src/VX_mem_coalescer.sv:178:5
	wire out_rsp_fire = out_rsp_valid && out_rsp_ready;
	// Trace: src/VX_mem_coalescer.sv:179:5
	wire out_rsp_eop;
	// Trace: src/VX_mem_coalescer.sv:180:5
	wire req_sent = state_r == STATE_SEND;
	// Trace: src/VX_mem_coalescer.sv:181:5
	assign ibuf_push = req_sent && ~in_req_rw;
	// Trace: src/VX_mem_coalescer.sv:182:5
	assign ibuf_pop = out_rsp_fire && out_rsp_eop;
	// Trace: src/VX_mem_coalescer.sv:183:5
	assign ibuf_raddr = out_rsp_tag[QUEUE_ADDRW - 1:0];
	// Trace: src/VX_mem_coalescer.sv:184:5
	wire [TAG_ID_WIDTH - 1:0] ibuf_din_tag = in_req_tag[TAG_ID_WIDTH - 1:0];
	// Trace: src/VX_mem_coalescer.sv:185:5
	wire [(NUM_REQS * DATA_RATIO_W) - 1:0] ibuf_din_offset = in_addr_offset;
	// Trace: src/VX_mem_coalescer.sv:186:5
	wire [NUM_REQS - 1:0] ibuf_din_pmask = current_pmask;
	// Trace: src/VX_mem_coalescer.sv:187:5
	assign ibuf_din = {ibuf_din_tag, ibuf_din_pmask, ibuf_din_offset};
	// Trace: src/VX_mem_coalescer.sv:188:5
	VX_index_buffer #(
		.DATAW(IBUF_DATA_WIDTH),
		.SIZE(QUEUE_SIZE)
	) req_ibuf(
		.clk(clk),
		.reset(reset),
		.acquire_en(ibuf_push),
		.write_addr(ibuf_waddr),
		.write_data(ibuf_din),
		.read_data(ibuf_dout),
		.read_addr(ibuf_raddr),
		.release_en(ibuf_pop),
		.full(ibuf_full),
		.empty(ibuf_empty)
	);
	// Trace: src/VX_mem_coalescer.sv:203:5
	assign out_req_valid = out_req_valid_r;
	// Trace: src/VX_mem_coalescer.sv:204:5
	assign out_req_rw = out_req_rw_r;
	// Trace: src/VX_mem_coalescer.sv:205:5
	assign out_req_mask = out_req_mask_r;
	// Trace: src/VX_mem_coalescer.sv:206:5
	assign out_req_byteen = out_req_byteen_r;
	// Trace: src/VX_mem_coalescer.sv:207:5
	assign out_req_addr = out_req_addr_r;
	// Trace: src/VX_mem_coalescer.sv:208:5
	generate
		if (FLAGS_WIDTH != 0) begin : g_out_req_flags
			// Trace: src/VX_mem_coalescer.sv:209:9
			assign out_req_flags = out_req_flags_r;
		end
		else begin : g_out_req_flags_0
			// Trace: src/VX_mem_coalescer.sv:211:9
			assign out_req_flags = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:213:5
	assign out_req_data = out_req_data_r;
	// Trace: src/VX_mem_coalescer.sv:214:5
	assign out_req_tag = out_req_tag_r;
	// Trace: src/VX_mem_coalescer.sv:215:5
	assign in_req_ready = in_req_ready_n;
	// Trace: src/VX_mem_coalescer.sv:216:5
	reg [(QUEUE_SIZE * OUT_REQS) - 1:0] rsp_rem_mask;
	// Trace: src/VX_mem_coalescer.sv:217:5
	wire [OUT_REQS - 1:0] rsp_rem_mask_n = rsp_rem_mask[ibuf_raddr * OUT_REQS+:OUT_REQS] & ~out_rsp_mask;
	// Trace: src/VX_mem_coalescer.sv:218:5
	assign out_rsp_eop = ~(|rsp_rem_mask_n);
	// Trace: src/VX_mem_coalescer.sv:219:5
	always @(posedge clk) begin
		// Trace: src/VX_mem_coalescer.sv:220:9
		if (ibuf_push)
			// Trace: src/VX_mem_coalescer.sv:221:13
			rsp_rem_mask[ibuf_waddr * OUT_REQS+:OUT_REQS] <= batch_valid_r;
		if (out_rsp_fire)
			// Trace: src/VX_mem_coalescer.sv:224:13
			rsp_rem_mask[ibuf_raddr * OUT_REQS+:OUT_REQS] <= rsp_rem_mask_n;
	end
	// Trace: src/VX_mem_coalescer.sv:227:5
	wire [(NUM_REQS * DATA_RATIO_W) - 1:0] ibuf_dout_offset;
	// Trace: src/VX_mem_coalescer.sv:228:5
	wire [NUM_REQS - 1:0] ibuf_dout_pmask;
	// Trace: src/VX_mem_coalescer.sv:229:5
	wire [TAG_ID_WIDTH - 1:0] ibuf_dout_tag;
	// Trace: src/VX_mem_coalescer.sv:230:5
	assign {ibuf_dout_tag, ibuf_dout_pmask, ibuf_dout_offset} = ibuf_dout;
	// Trace: src/VX_mem_coalescer.sv:231:5
	wire [(NUM_REQS * DATA_IN_WIDTH) - 1:0] in_rsp_data_n;
	// Trace: src/VX_mem_coalescer.sv:232:5
	genvar _gv_i_104;
	generate
		for (_gv_i_104 = 0; _gv_i_104 < OUT_REQS; _gv_i_104 = _gv_i_104 + 1) begin : g_in_rsp_data_n
			localparam i = _gv_i_104;
			genvar _gv_j_14;
			for (_gv_j_14 = 0; _gv_j_14 < DATA_RATIO; _gv_j_14 = _gv_j_14 + 1) begin : g_j
				localparam j = _gv_j_14;
				// Trace: src/VX_mem_coalescer.sv:234:13
				assign in_rsp_data_n[((i * DATA_RATIO) + j) * DATA_IN_WIDTH+:DATA_IN_WIDTH] = out_rsp_data[(i * DATA_OUT_WIDTH) + (ibuf_dout_offset[((i * DATA_RATIO) + j) * DATA_RATIO_W+:DATA_RATIO_W] * DATA_IN_WIDTH)+:DATA_IN_WIDTH];
			end
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:237:5
	wire [NUM_REQS - 1:0] in_rsp_mask_n;
	// Trace: src/VX_mem_coalescer.sv:238:5
	genvar _gv_i_105;
	generate
		for (_gv_i_105 = 0; _gv_i_105 < OUT_REQS; _gv_i_105 = _gv_i_105 + 1) begin : g_in_rsp_mask_n
			localparam i = _gv_i_105;
			genvar _gv_j_15;
			for (_gv_j_15 = 0; _gv_j_15 < DATA_RATIO; _gv_j_15 = _gv_j_15 + 1) begin : g_j
				localparam j = _gv_j_15;
				// Trace: src/VX_mem_coalescer.sv:240:13
				assign in_rsp_mask_n[(i * DATA_RATIO) + j] = out_rsp_mask[i] && ibuf_dout_pmask[(i * DATA_RATIO) + j];
			end
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:243:5
	assign in_rsp_valid = out_rsp_valid;
	// Trace: src/VX_mem_coalescer.sv:244:5
	assign in_rsp_mask = in_rsp_mask_n;
	// Trace: src/VX_mem_coalescer.sv:245:5
	assign in_rsp_data = in_rsp_data_n;
	// Trace: src/VX_mem_coalescer.sv:246:5
	assign in_rsp_tag = {out_rsp_tag[OUT_TAG_WIDTH - 1-:UUID_WIDTH], ibuf_dout_tag};
	// Trace: src/VX_mem_coalescer.sv:247:5
	assign out_rsp_ready = in_rsp_ready;
endmodule
module VX_stream_pack (
	clk,
	reset,
	valid_in,
	data_in,
	tag_in,
	ready_in,
	valid_out,
	mask_out,
	data_out,
	tag_out,
	ready_out
);
	// Trace: src/VX_stream_pack.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_stream_pack.sv:3:15
	parameter DATA_WIDTH = 1;
	// Trace: src/VX_stream_pack.sv:4:15
	parameter TAG_WIDTH = 1;
	// Trace: src/VX_stream_pack.sv:5:15
	parameter TAG_SEL_BITS = 0;
	// Trace: src/VX_stream_pack.sv:6:15
	parameter ARBITER = "P";
	// Trace: src/VX_stream_pack.sv:7:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_pack.sv:9:5
	input wire clk;
	// Trace: src/VX_stream_pack.sv:10:5
	input wire reset;
	// Trace: src/VX_stream_pack.sv:11:5
	input wire [NUM_REQS - 1:0] valid_in;
	// Trace: src/VX_stream_pack.sv:12:5
	input wire [(NUM_REQS * DATA_WIDTH) - 1:0] data_in;
	// Trace: src/VX_stream_pack.sv:13:5
	input wire [(NUM_REQS * TAG_WIDTH) - 1:0] tag_in;
	// Trace: src/VX_stream_pack.sv:14:5
	output wire [NUM_REQS - 1:0] ready_in;
	// Trace: src/VX_stream_pack.sv:15:5
	output wire valid_out;
	// Trace: src/VX_stream_pack.sv:16:5
	output wire [NUM_REQS - 1:0] mask_out;
	// Trace: src/VX_stream_pack.sv:17:5
	output wire [(NUM_REQS * DATA_WIDTH) - 1:0] data_out;
	// Trace: src/VX_stream_pack.sv:18:5
	output wire [TAG_WIDTH - 1:0] tag_out;
	// Trace: src/VX_stream_pack.sv:19:5
	input wire ready_out;
	// Trace: src/VX_stream_pack.sv:21:5
	generate
		if (NUM_REQS > 1) begin : g_pack
			// Trace: src/VX_stream_pack.sv:22:9
			localparam LOG_NUM_REQS = $clog2(NUM_REQS);
			// Trace: src/VX_stream_pack.sv:23:9
			wire [LOG_NUM_REQS - 1:0] grant_index;
			// Trace: src/VX_stream_pack.sv:24:9
			wire grant_valid;
			// Trace: src/VX_stream_pack.sv:25:9
			wire grant_ready;
			// Trace: src/VX_stream_pack.sv:26:9
			VX_generic_arbiter #(
				.NUM_REQS(NUM_REQS),
				.TYPE(ARBITER)
			) arbiter(
				.clk(clk),
				.reset(reset),
				.requests(valid_in),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(),
				.grant_ready(grant_ready)
			);
			// Trace: src/VX_stream_pack.sv:38:9
			wire [TAG_WIDTH - 1:0] tag_sel = tag_in[grant_index * TAG_WIDTH+:TAG_WIDTH];
			// Trace: src/VX_stream_pack.sv:39:9
			wire [NUM_REQS - 1:0] tag_matches;
			genvar _gv_i_106;
			for (_gv_i_106 = 0; _gv_i_106 < NUM_REQS; _gv_i_106 = _gv_i_106 + 1) begin : g_tag_matches
				localparam i = _gv_i_106;
				// Trace: src/VX_stream_pack.sv:41:13
				assign tag_matches[i] = tag_in[(i * TAG_WIDTH) + (TAG_SEL_BITS - 1)-:TAG_SEL_BITS] == tag_sel[TAG_SEL_BITS - 1:0];
			end
			genvar _gv_i_107;
			for (_gv_i_107 = 0; _gv_i_107 < NUM_REQS; _gv_i_107 = _gv_i_107 + 1) begin : g_ready_in
				localparam i = _gv_i_107;
				// Trace: src/VX_stream_pack.sv:44:13
				assign ready_in[i] = grant_ready & tag_matches[i];
			end
			// Trace: src/VX_stream_pack.sv:46:9
			wire [NUM_REQS - 1:0] mask_sel = valid_in & tag_matches;
			// Trace: src/VX_stream_pack.sv:47:9
			VX_elastic_buffer #(
				.DATAW((NUM_REQS + TAG_WIDTH) + (NUM_REQS * DATA_WIDTH)),
				.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
				.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
			) out_buf(
				.clk(clk),
				.reset(reset),
				.valid_in(grant_valid),
				.data_in({mask_sel, tag_sel, data_in}),
				.ready_in(grant_ready),
				.valid_out(valid_out),
				.data_out({mask_out, tag_out, data_out}),
				.ready_out(ready_out)
			);
		end
		else begin : g_passthru
			// Trace: src/VX_stream_pack.sv:62:9
			assign valid_out = valid_in;
			// Trace: src/VX_stream_pack.sv:63:9
			assign mask_out = 1'b1;
			// Trace: src/VX_stream_pack.sv:64:9
			assign data_out = data_in;
			// Trace: src/VX_stream_pack.sv:65:9
			assign tag_out = tag_in;
			// Trace: src/VX_stream_pack.sv:66:9
			assign ready_in = ready_out;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_cache_flush
module VX_cache_tags (
	clk,
	reset,
	init,
	flush,
	fill,
	read,
	write,
	line_idx,
	line_tag,
	evict_way,
	tag_matches,
	evict_dirty,
	evict_tag
);
	// Trace: src/VX_cache_tags.sv:2:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_cache_tags.sv:3:15
	parameter LINE_SIZE = 16;
	// Trace: src/VX_cache_tags.sv:4:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_tags.sv:5:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_tags.sv:6:15
	parameter WORD_SIZE = 1;
	// Trace: src/VX_cache_tags.sv:7:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_cache_tags.sv:9:5
	input wire clk;
	// Trace: src/VX_cache_tags.sv:10:5
	input wire reset;
	// Trace: src/VX_cache_tags.sv:11:5
	input wire init;
	// Trace: src/VX_cache_tags.sv:12:5
	input wire flush;
	// Trace: src/VX_cache_tags.sv:13:5
	input wire fill;
	// Trace: src/VX_cache_tags.sv:14:5
	input wire read;
	// Trace: src/VX_cache_tags.sv:15:5
	input wire write;
	// Trace: src/VX_cache_tags.sv:16:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx;
	// Trace: src/VX_cache_tags.sv:17:5
	input wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] line_tag;
	// Trace: src/VX_cache_tags.sv:18:5
	input wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] evict_way;
	// Trace: src/VX_cache_tags.sv:19:5
	output wire [NUM_WAYS - 1:0] tag_matches;
	// Trace: src/VX_cache_tags.sv:20:5
	output wire evict_dirty;
	// Trace: src/VX_cache_tags.sv:21:5
	output wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] evict_tag;
	// Trace: src/VX_cache_tags.sv:23:5
	localparam TAG_WIDTH = (1 + WRITEBACK) + (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1));
	// Trace: src/VX_cache_tags.sv:24:5
	wire [(NUM_WAYS * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))) - 1:0] read_tag;
	// Trace: src/VX_cache_tags.sv:25:5
	wire [NUM_WAYS - 1:0] read_valid;
	// Trace: src/VX_cache_tags.sv:26:5
	wire [NUM_WAYS - 1:0] read_dirty;
	// Trace: src/VX_cache_tags.sv:27:5
	generate
		if (WRITEBACK) begin : g_evict_tag_wb
			// Trace: src/VX_cache_tags.sv:28:9
			assign evict_dirty = read_dirty[evict_way];
			// Trace: src/VX_cache_tags.sv:29:9
			assign evict_tag = read_tag[evict_way * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))+:((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)];
		end
		else begin : g_evict_tag_wt
			// Trace: src/VX_cache_tags.sv:31:9
			assign evict_dirty = 1'b0;
			// Trace: src/VX_cache_tags.sv:32:9
			assign evict_tag = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_cache_tags.sv:34:5
	genvar _gv_i_121;
	generate
		for (_gv_i_121 = 0; _gv_i_121 < NUM_WAYS; _gv_i_121 = _gv_i_121 + 1) begin : g_tag_store
			localparam i = _gv_i_121;
			// Trace: src/VX_cache_tags.sv:35:9
			wire way_en = (NUM_WAYS == 1) || (evict_way == i);
			// Trace: src/VX_cache_tags.sv:36:9
			wire do_init = init;
			// Trace: src/VX_cache_tags.sv:37:9
			wire do_fill = fill && way_en;
			// Trace: src/VX_cache_tags.sv:38:9
			wire do_flush = flush && (!WRITEBACK || way_en);
			// Trace: src/VX_cache_tags.sv:39:9
			wire do_write = (WRITEBACK && write) && tag_matches[i];
			// Trace: src/VX_cache_tags.sv:40:9
			wire line_read = (read || write) || (WRITEBACK && (fill || flush));
			// Trace: src/VX_cache_tags.sv:41:9
			wire line_write = ((do_init || do_fill) || do_flush) || do_write;
			// Trace: src/VX_cache_tags.sv:42:9
			wire line_valid = fill || write;
			// Trace: src/VX_cache_tags.sv:43:9
			wire [TAG_WIDTH - 1:0] line_wdata;
			// Trace: src/VX_cache_tags.sv:44:9
			wire [TAG_WIDTH - 1:0] line_rdata;
			if (WRITEBACK) begin : g_wdata
				// Trace: src/VX_cache_tags.sv:46:13
				assign line_wdata = {line_valid, write, line_tag};
				// Trace: src/VX_cache_tags.sv:47:13
				assign {read_valid[i], read_dirty[i], read_tag[i * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))+:((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)]} = line_rdata;
			end
			else begin : g_wdata
				// Trace: src/VX_cache_tags.sv:49:13
				assign line_wdata = {line_valid, line_tag};
				// Trace: src/VX_cache_tags.sv:50:13
				assign {read_valid[i], read_tag[i * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))+:((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)]} = line_rdata;
				// Trace: src/VX_cache_tags.sv:51:13
				assign read_dirty[i] = 1'b0;
			end
			// Trace: src/VX_cache_tags.sv:53:9
			VX_sp_ram #(
				.DATAW(TAG_WIDTH),
				.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
				.RDW_MODE("W"),
				.RADDR_REG(1)
			) tag_store(
				.clk(clk),
				.reset(reset),
				.read(line_read),
				.write(line_write),
				.wren(1'b1),
				.addr(line_idx),
				.wdata(line_wdata),
				.rdata(line_rdata)
			);
		end
	endgenerate
	// Trace: src/VX_cache_tags.sv:69:5
	genvar _gv_i_122;
	generate
		for (_gv_i_122 = 0; _gv_i_122 < NUM_WAYS; _gv_i_122 = _gv_i_122 + 1) begin : g_tag_matches
			localparam i = _gv_i_122;
			// Trace: src/VX_cache_tags.sv:70:9
			assign tag_matches[i] = read_valid[i] && (line_tag == read_tag[i * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))+:((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)]);
		end
	endgenerate
endmodule
// removed interface: VX_warp_ctl_if
module Vortex (
	clk,
	reset,
	mem_req_valid,
	mem_req_rw,
	mem_req_byteen,
	mem_req_addr,
	mem_req_data,
	mem_req_tag,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready,
	dcr_wr_valid,
	dcr_wr_addr,
	dcr_wr_data,
	busy
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/Vortex.sv:2:5
	input wire clk;
	// Trace: src/Vortex.sv:3:5
	input wire reset;
	// Trace: src/Vortex.sv:4:5
	localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
	localparam VX_gpu_pkg_LSU_WORD_SIZE = 4;
	localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
	localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
	localparam VX_gpu_pkg_L2_NUM_REQS = 1;
	localparam VX_gpu_pkg_L3_NUM_REQS = 1;
	output wire [0:0] mem_req_valid;
	// Trace: src/Vortex.sv:5:5
	output wire [0:0] mem_req_rw;
	// Trace: src/Vortex.sv:6:5
	output wire [63:0] mem_req_byteen;
	// Trace: src/Vortex.sv:7:5
	output wire [25:0] mem_req_addr;
	// Trace: src/Vortex.sv:8:5
	output wire [511:0] mem_req_data;
	// Trace: src/Vortex.sv:9:5
	localparam VX_gpu_pkg_DCACHE_LINE_SIZE = 64;
	localparam VX_gpu_pkg_DCACHE_MERGED_REQS = 1;
	localparam VX_gpu_pkg_DCACHE_MEM_BATCHES = 1;
	localparam VX_gpu_pkg_DCACHE_TAG_ID_BITS = 2;
	localparam VX_gpu_pkg_DCACHE_TAG_WIDTH = 3;
	localparam VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH = 6;
	localparam VX_gpu_pkg_ICACHE_MEM_TAG_WIDTH = 5;
	localparam VX_gpu_pkg_L1_MEM_TAG_WIDTH = VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH;
	localparam VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH = 7;
	localparam VX_gpu_pkg_L2_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
	localparam VX_gpu_pkg_L2_WORD_SIZE = 64;
	localparam VX_gpu_pkg_L2_MEM_TAG_WIDTH = 7;
	localparam VX_gpu_pkg_L3_TAG_WIDTH = VX_gpu_pkg_L2_MEM_TAG_WIDTH;
	localparam VX_gpu_pkg_L3_WORD_SIZE = 64;
	localparam VX_gpu_pkg_L3_MEM_TAG_WIDTH = 7;
	output wire [6:0] mem_req_tag;
	// Trace: src/Vortex.sv:10:5
	input wire [0:0] mem_req_ready;
	// Trace: src/Vortex.sv:11:5
	input wire [0:0] mem_rsp_valid;
	// Trace: src/Vortex.sv:12:5
	input wire [511:0] mem_rsp_data;
	// Trace: src/Vortex.sv:13:5
	input wire [6:0] mem_rsp_tag;
	// Trace: src/Vortex.sv:14:5
	output wire [0:0] mem_rsp_ready;
	// Trace: src/Vortex.sv:15:5
	input wire dcr_wr_valid;
	// Trace: src/Vortex.sv:16:5
	input wire [11:0] dcr_wr_addr;
	// Trace: src/Vortex.sv:17:5
	input wire [31:0] dcr_wr_data;
	// Trace: src/Vortex.sv:18:5
	output wire busy;
	// Trace: src/Vortex.sv:20:5
	// expanded interface instance: per_cluster_mem_bus_if
	localparam _param_CA4E3_DATA_SIZE = 64;
	localparam _param_CA4E3_TAG_WIDTH = VX_gpu_pkg_L2_MEM_TAG_WIDTH;
	genvar _arr_CA4E3;
	generate
		for (_arr_CA4E3 = 0; _arr_CA4E3 <= 0; _arr_CA4E3 = _arr_CA4E3 + 1) begin : per_cluster_mem_bus_if
			// Trace: src/VX_mem_bus_if.sv:2:15
			localparam DATA_SIZE = _param_CA4E3_DATA_SIZE;
			// Trace: src/VX_mem_bus_if.sv:3:15
			localparam FLAGS_WIDTH = 3;
			// Trace: src/VX_mem_bus_if.sv:4:15
			localparam TAG_WIDTH = _param_CA4E3_TAG_WIDTH;
			// Trace: src/VX_mem_bus_if.sv:5:15
			localparam MEM_ADDR_WIDTH = 32;
			// Trace: src/VX_mem_bus_if.sv:6:15
			localparam ADDR_WIDTH = 26;
			// Trace: src/VX_mem_bus_if.sv:7:15
			localparam UUID_WIDTH = 1;
			// Trace: src/VX_mem_bus_if.sv:9:5
			// removed localparam type tag_t
			// Trace: src/VX_mem_bus_if.sv:13:5
			// removed localparam type req_data_t
			// Trace: src/VX_mem_bus_if.sv:21:5
			// removed localparam type rsp_data_t
			// Trace: src/VX_mem_bus_if.sv:25:5
			wire req_valid;
			// Trace: src/VX_mem_bus_if.sv:26:5
			wire [612:0] req_data;
			// Trace: src/VX_mem_bus_if.sv:27:5
			wire req_ready;
			// Trace: src/VX_mem_bus_if.sv:28:5
			wire rsp_valid;
			// Trace: src/VX_mem_bus_if.sv:29:5
			wire [518:0] rsp_data;
			// Trace: src/VX_mem_bus_if.sv:30:5
			wire rsp_ready;
			// Trace: src/VX_mem_bus_if.sv:31:5
			// Trace: src/VX_mem_bus_if.sv:39:5
		end
	endgenerate
	// Trace: src/Vortex.sv:24:5
	// expanded interface instance: mem_bus_if
	localparam _param_4F26C_DATA_SIZE = 64;
	localparam _param_4F26C_TAG_WIDTH = VX_gpu_pkg_L3_MEM_TAG_WIDTH;
	genvar _arr_4F26C;
	generate
		for (_arr_4F26C = 0; _arr_4F26C <= 0; _arr_4F26C = _arr_4F26C + 1) begin : mem_bus_if
			// Trace: src/VX_mem_bus_if.sv:2:15
			localparam DATA_SIZE = _param_4F26C_DATA_SIZE;
			// Trace: src/VX_mem_bus_if.sv:3:15
			localparam FLAGS_WIDTH = 3;
			// Trace: src/VX_mem_bus_if.sv:4:15
			localparam TAG_WIDTH = _param_4F26C_TAG_WIDTH;
			// Trace: src/VX_mem_bus_if.sv:5:15
			localparam MEM_ADDR_WIDTH = 32;
			// Trace: src/VX_mem_bus_if.sv:6:15
			localparam ADDR_WIDTH = 26;
			// Trace: src/VX_mem_bus_if.sv:7:15
			localparam UUID_WIDTH = 1;
			// Trace: src/VX_mem_bus_if.sv:9:5
			// removed localparam type tag_t
			// Trace: src/VX_mem_bus_if.sv:13:5
			// removed localparam type req_data_t
			// Trace: src/VX_mem_bus_if.sv:21:5
			// removed localparam type rsp_data_t
			// Trace: src/VX_mem_bus_if.sv:25:5
			wire req_valid;
			// Trace: src/VX_mem_bus_if.sv:26:5
			wire [612:0] req_data;
			// Trace: src/VX_mem_bus_if.sv:27:5
			wire req_ready;
			// Trace: src/VX_mem_bus_if.sv:28:5
			wire rsp_valid;
			// Trace: src/VX_mem_bus_if.sv:29:5
			wire [518:0] rsp_data;
			// Trace: src/VX_mem_bus_if.sv:30:5
			wire rsp_ready;
			// Trace: src/VX_mem_bus_if.sv:31:5
			// Trace: src/VX_mem_bus_if.sv:39:5
		end
	endgenerate
	// Trace: src/Vortex.sv:28:5
	wire [0:0] l3_reset;
	// Trace: src/Vortex.sv:29:5
	VX_reset_relay #(
		.N(1),
		.MAX_FANOUT(0)
	) __l3_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(l3_reset)
	);
	// Trace: src/Vortex.sv:34:5
	// expanded module instance: l3cache
	localparam _bbase_56375_core_bus_if = 0;
	localparam _bbase_56375_mem_bus_if = 0;
	localparam _param_56375_INSTANCE_ID = "l3cache";
	localparam _param_56375_CACHE_SIZE = 2097152;
	localparam _param_56375_LINE_SIZE = 64;
	localparam _param_56375_NUM_BANKS = VX_gpu_pkg_L3_NUM_REQS;
	localparam _param_56375_NUM_WAYS = 8;
	localparam _param_56375_WORD_SIZE = VX_gpu_pkg_L3_WORD_SIZE;
	localparam _param_56375_NUM_REQS = VX_gpu_pkg_L3_NUM_REQS;
	localparam _param_56375_MEM_PORTS = VX_gpu_pkg_L3_NUM_REQS;
	localparam _param_56375_CRSQ_SIZE = 2;
	localparam _param_56375_MSHR_SIZE = 16;
	localparam _param_56375_MRSQ_SIZE = 4;
	localparam _param_56375_MREQ_SIZE = 4;
	localparam _param_56375_TAG_WIDTH = VX_gpu_pkg_L2_MEM_TAG_WIDTH;
	localparam _param_56375_WRITE_ENABLE = 1;
	localparam _param_56375_WRITEBACK = 0;
	localparam _param_56375_DIRTY_BYTES = 0;
	localparam _param_56375_REPL_POLICY = 1;
	localparam _param_56375_UUID_WIDTH = 1;
	localparam _param_56375_FLAGS_WIDTH = 3;
	localparam _param_56375_CORE_OUT_BUF = 3;
	localparam _param_56375_MEM_OUT_BUF = 3;
	localparam _param_56375_NC_ENABLE = 1;
	localparam _param_56375_PASSTHRU = 1'd1;
	function automatic [6:0] sv2v_cast_7;
		input reg [6:0] inp;
		sv2v_cast_7 = inp;
	endfunction
	generate
		if (1) begin : l3cache
			// removed import VX_gpu_pkg::*;
			// Trace: src/VX_cache_wrap.sv:2:16
			localparam INSTANCE_ID = _param_56375_INSTANCE_ID;
			// Trace: src/VX_cache_wrap.sv:3:15
			localparam TAG_SEL_IDX = 0;
			// Trace: src/VX_cache_wrap.sv:4:15
			localparam NUM_REQS = _param_56375_NUM_REQS;
			// Trace: src/VX_cache_wrap.sv:5:15
			localparam MEM_PORTS = _param_56375_MEM_PORTS;
			// Trace: src/VX_cache_wrap.sv:6:15
			localparam CACHE_SIZE = _param_56375_CACHE_SIZE;
			// Trace: src/VX_cache_wrap.sv:7:15
			localparam LINE_SIZE = _param_56375_LINE_SIZE;
			// Trace: src/VX_cache_wrap.sv:8:15
			localparam NUM_BANKS = _param_56375_NUM_BANKS;
			// Trace: src/VX_cache_wrap.sv:9:15
			localparam NUM_WAYS = _param_56375_NUM_WAYS;
			// Trace: src/VX_cache_wrap.sv:10:15
			localparam WORD_SIZE = _param_56375_WORD_SIZE;
			// Trace: src/VX_cache_wrap.sv:11:15
			localparam CRSQ_SIZE = _param_56375_CRSQ_SIZE;
			// Trace: src/VX_cache_wrap.sv:12:15
			localparam MSHR_SIZE = _param_56375_MSHR_SIZE;
			// Trace: src/VX_cache_wrap.sv:13:15
			localparam MRSQ_SIZE = _param_56375_MRSQ_SIZE;
			// Trace: src/VX_cache_wrap.sv:14:15
			localparam MREQ_SIZE = _param_56375_MREQ_SIZE;
			// Trace: src/VX_cache_wrap.sv:15:15
			localparam WRITE_ENABLE = _param_56375_WRITE_ENABLE;
			// Trace: src/VX_cache_wrap.sv:16:15
			localparam WRITEBACK = _param_56375_WRITEBACK;
			// Trace: src/VX_cache_wrap.sv:17:15
			localparam DIRTY_BYTES = _param_56375_DIRTY_BYTES;
			// Trace: src/VX_cache_wrap.sv:18:15
			localparam REPL_POLICY = _param_56375_REPL_POLICY;
			// Trace: src/VX_cache_wrap.sv:19:15
			localparam UUID_WIDTH = _param_56375_UUID_WIDTH;
			// Trace: src/VX_cache_wrap.sv:20:15
			localparam TAG_WIDTH = _param_56375_TAG_WIDTH;
			// Trace: src/VX_cache_wrap.sv:21:15
			localparam FLAGS_WIDTH = _param_56375_FLAGS_WIDTH;
			// Trace: src/VX_cache_wrap.sv:22:15
			localparam NC_ENABLE = _param_56375_NC_ENABLE;
			// Trace: src/VX_cache_wrap.sv:23:15
			localparam PASSTHRU = _param_56375_PASSTHRU;
			// Trace: src/VX_cache_wrap.sv:24:15
			localparam CORE_OUT_BUF = _param_56375_CORE_OUT_BUF;
			// Trace: src/VX_cache_wrap.sv:25:15
			localparam MEM_OUT_BUF = _param_56375_MEM_OUT_BUF;
			// Trace: src/VX_cache_wrap.sv:27:5
			wire clk;
			// Trace: src/VX_cache_wrap.sv:28:5
			wire reset;
			// Trace: src/VX_cache_wrap.sv:29:5
			localparam _mbase_core_bus_if = 0;
			// Trace: src/VX_cache_wrap.sv:30:5
			localparam _mbase_mem_bus_if = 0;
			// Trace: src/VX_cache_wrap.sv:32:5
			localparam CACHE_MEM_TAG_WIDTH = 5;
			// Trace: src/VX_cache_wrap.sv:34:5
			localparam BYPASS_TAG_WIDTH = 7;
			// Trace: src/VX_cache_wrap.sv:36:5
			localparam NC_TAG_WIDTH = 8;
			// Trace: src/VX_cache_wrap.sv:37:5
			localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
			// Trace: src/VX_cache_wrap.sv:38:5
			localparam BYPASS_ENABLE = 1'd1;
			// Trace: src/VX_cache_wrap.sv:39:5
			// expanded interface instance: core_bus_cache_if
			localparam _param_24C1C_DATA_SIZE = WORD_SIZE;
			localparam _param_24C1C_TAG_WIDTH = TAG_WIDTH;
			genvar _arr_24C1C;
			for (_arr_24C1C = 0; _arr_24C1C <= 0; _arr_24C1C = _arr_24C1C + 1) begin : core_bus_cache_if
				// Trace: src/VX_mem_bus_if.sv:2:15
				localparam DATA_SIZE = _param_24C1C_DATA_SIZE;
				// Trace: src/VX_mem_bus_if.sv:3:15
				localparam FLAGS_WIDTH = 3;
				// Trace: src/VX_mem_bus_if.sv:4:15
				localparam TAG_WIDTH = _param_24C1C_TAG_WIDTH;
				// Trace: src/VX_mem_bus_if.sv:5:15
				localparam MEM_ADDR_WIDTH = 32;
				// Trace: src/VX_mem_bus_if.sv:6:15
				localparam ADDR_WIDTH = 26;
				// Trace: src/VX_mem_bus_if.sv:7:15
				localparam UUID_WIDTH = 1;
				// Trace: src/VX_mem_bus_if.sv:9:5
				// removed localparam type tag_t
				// Trace: src/VX_mem_bus_if.sv:13:5
				// removed localparam type req_data_t
				// Trace: src/VX_mem_bus_if.sv:21:5
				// removed localparam type rsp_data_t
				// Trace: src/VX_mem_bus_if.sv:25:5
				wire req_valid;
				// Trace: src/VX_mem_bus_if.sv:26:5
				wire [612:0] req_data;
				// Trace: src/VX_mem_bus_if.sv:27:5
				wire req_ready;
				// Trace: src/VX_mem_bus_if.sv:28:5
				wire rsp_valid;
				// Trace: src/VX_mem_bus_if.sv:29:5
				wire [518:0] rsp_data;
				// Trace: src/VX_mem_bus_if.sv:30:5
				wire rsp_ready;
				// Trace: src/VX_mem_bus_if.sv:31:5
				// Trace: src/VX_mem_bus_if.sv:39:5
			end
			// Trace: src/VX_cache_wrap.sv:43:5
			// expanded interface instance: mem_bus_cache_if
			localparam _param_D895D_DATA_SIZE = LINE_SIZE;
			localparam _param_D895D_TAG_WIDTH = CACHE_MEM_TAG_WIDTH;
			genvar _arr_D895D;
			for (_arr_D895D = 0; _arr_D895D <= 0; _arr_D895D = _arr_D895D + 1) begin : mem_bus_cache_if
				// Trace: src/VX_mem_bus_if.sv:2:15
				localparam DATA_SIZE = _param_D895D_DATA_SIZE;
				// Trace: src/VX_mem_bus_if.sv:3:15
				localparam FLAGS_WIDTH = 3;
				// Trace: src/VX_mem_bus_if.sv:4:15
				localparam TAG_WIDTH = _param_D895D_TAG_WIDTH;
				// Trace: src/VX_mem_bus_if.sv:5:15
				localparam MEM_ADDR_WIDTH = 32;
				// Trace: src/VX_mem_bus_if.sv:6:15
				localparam ADDR_WIDTH = 26;
				// Trace: src/VX_mem_bus_if.sv:7:15
				localparam UUID_WIDTH = 1;
				// Trace: src/VX_mem_bus_if.sv:9:5
				// removed localparam type tag_t
				// Trace: src/VX_mem_bus_if.sv:13:5
				// removed localparam type req_data_t
				// Trace: src/VX_mem_bus_if.sv:21:5
				// removed localparam type rsp_data_t
				// Trace: src/VX_mem_bus_if.sv:25:5
				wire req_valid;
				// Trace: src/VX_mem_bus_if.sv:26:5
				wire [610:0] req_data;
				// Trace: src/VX_mem_bus_if.sv:27:5
				wire req_ready;
				// Trace: src/VX_mem_bus_if.sv:28:5
				wire rsp_valid;
				// Trace: src/VX_mem_bus_if.sv:29:5
				wire [516:0] rsp_data;
				// Trace: src/VX_mem_bus_if.sv:30:5
				wire rsp_ready;
				// Trace: src/VX_mem_bus_if.sv:31:5
				// Trace: src/VX_mem_bus_if.sv:39:5
			end
			// Trace: src/VX_cache_wrap.sv:47:5
			// expanded interface instance: mem_bus_tmp_if
			localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
			localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
			genvar _arr_4FE36;
			for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
				// Trace: src/VX_mem_bus_if.sv:2:15
				localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
				// Trace: src/VX_mem_bus_if.sv:3:15
				localparam FLAGS_WIDTH = 3;
				// Trace: src/VX_mem_bus_if.sv:4:15
				localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
				// Trace: src/VX_mem_bus_if.sv:5:15
				localparam MEM_ADDR_WIDTH = 32;
				// Trace: src/VX_mem_bus_if.sv:6:15
				localparam ADDR_WIDTH = 26;
				// Trace: src/VX_mem_bus_if.sv:7:15
				localparam UUID_WIDTH = 1;
				// Trace: src/VX_mem_bus_if.sv:9:5
				// removed localparam type tag_t
				// Trace: src/VX_mem_bus_if.sv:13:5
				// removed localparam type req_data_t
				// Trace: src/VX_mem_bus_if.sv:21:5
				// removed localparam type rsp_data_t
				// Trace: src/VX_mem_bus_if.sv:25:5
				wire req_valid;
				// Trace: src/VX_mem_bus_if.sv:26:5
				wire [(606 + (_param_4FE36_TAG_WIDTH + 0)) - 1:0] req_data;
				// Trace: src/VX_mem_bus_if.sv:27:5
				wire req_ready;
				// Trace: src/VX_mem_bus_if.sv:28:5
				wire rsp_valid;
				// Trace: src/VX_mem_bus_if.sv:29:5
				wire [(512 + (_param_4FE36_TAG_WIDTH + 0)) - 1:0] rsp_data;
				// Trace: src/VX_mem_bus_if.sv:30:5
				wire rsp_ready;
				// Trace: src/VX_mem_bus_if.sv:31:5
				// Trace: src/VX_mem_bus_if.sv:39:5
			end
			// Trace: src/VX_cache_wrap.sv:51:5
			if (BYPASS_ENABLE) begin : g_bypass
				// Trace: src/VX_cache_wrap.sv:52:9
				// expanded module instance: cache_bypass
				localparam _bbase_714AA_core_bus_in_if = 0;
				localparam _bbase_714AA_core_bus_out_if = 0;
				localparam _bbase_714AA_mem_bus_in_if = 0;
				localparam _bbase_714AA_mem_bus_out_if = 0;
				localparam _param_714AA_NUM_REQS = NUM_REQS;
				localparam _param_714AA_MEM_PORTS = MEM_PORTS;
				localparam _param_714AA_TAG_SEL_IDX = TAG_SEL_IDX;
				localparam _param_714AA_CACHE_ENABLE = !PASSTHRU;
				localparam _param_714AA_WORD_SIZE = WORD_SIZE;
				localparam _param_714AA_LINE_SIZE = LINE_SIZE;
				localparam _param_714AA_CORE_ADDR_WIDTH = 26;
				localparam _param_714AA_CORE_TAG_WIDTH = TAG_WIDTH;
				localparam _param_714AA_MEM_ADDR_WIDTH = 26;
				localparam _param_714AA_MEM_TAG_IN_WIDTH = CACHE_MEM_TAG_WIDTH;
				localparam _param_714AA_UUID_WIDTH = UUID_WIDTH;
				localparam _param_714AA_CORE_OUT_BUF = CORE_OUT_BUF;
				localparam _param_714AA_MEM_OUT_BUF = MEM_OUT_BUF;
				if (1) begin : cache_bypass
					// Trace: src/VX_cache_bypass.sv:2:15
					localparam NUM_REQS = _param_714AA_NUM_REQS;
					// Trace: src/VX_cache_bypass.sv:3:15
					localparam MEM_PORTS = _param_714AA_MEM_PORTS;
					// Trace: src/VX_cache_bypass.sv:4:15
					localparam TAG_SEL_IDX = _param_714AA_TAG_SEL_IDX;
					// Trace: src/VX_cache_bypass.sv:5:15
					localparam CACHE_ENABLE = _param_714AA_CACHE_ENABLE;
					// Trace: src/VX_cache_bypass.sv:6:15
					localparam WORD_SIZE = _param_714AA_WORD_SIZE;
					// Trace: src/VX_cache_bypass.sv:7:15
					localparam LINE_SIZE = _param_714AA_LINE_SIZE;
					// Trace: src/VX_cache_bypass.sv:8:15
					localparam CORE_ADDR_WIDTH = _param_714AA_CORE_ADDR_WIDTH;
					// Trace: src/VX_cache_bypass.sv:9:15
					localparam CORE_TAG_WIDTH = _param_714AA_CORE_TAG_WIDTH;
					// Trace: src/VX_cache_bypass.sv:10:15
					localparam MEM_ADDR_WIDTH = _param_714AA_MEM_ADDR_WIDTH;
					// Trace: src/VX_cache_bypass.sv:11:15
					localparam MEM_TAG_IN_WIDTH = _param_714AA_MEM_TAG_IN_WIDTH;
					// Trace: src/VX_cache_bypass.sv:12:15
					localparam UUID_WIDTH = _param_714AA_UUID_WIDTH;
					// Trace: src/VX_cache_bypass.sv:13:15
					localparam CORE_OUT_BUF = _param_714AA_CORE_OUT_BUF;
					// Trace: src/VX_cache_bypass.sv:14:15
					localparam MEM_OUT_BUF = _param_714AA_MEM_OUT_BUF;
					// Trace: src/VX_cache_bypass.sv:16:5
					wire clk;
					// Trace: src/VX_cache_bypass.sv:17:5
					wire reset;
					// Trace: src/VX_cache_bypass.sv:18:5
					localparam _mbase_core_bus_in_if = 0;
					// Trace: src/VX_cache_bypass.sv:19:5
					localparam _mbase_core_bus_out_if = 0;
					// Trace: src/VX_cache_bypass.sv:20:5
					localparam _mbase_mem_bus_in_if = 0;
					// Trace: src/VX_cache_bypass.sv:21:5
					localparam _mbase_mem_bus_out_if = 0;
					// Trace: src/VX_cache_bypass.sv:23:5
					localparam DIRECT_PASSTHRU = (!CACHE_ENABLE && 1'd1) && 1'd1;
					// Trace: src/VX_cache_bypass.sv:24:5
					localparam CORE_DATA_WIDTH = 512;
					// Trace: src/VX_cache_bypass.sv:25:5
					localparam WORDS_PER_LINE = 1;
					// Trace: src/VX_cache_bypass.sv:26:5
					localparam WSEL_BITS = 0;
					// Trace: src/VX_cache_bypass.sv:27:5
					localparam CORE_TAG_ID_WIDTH = 6;
					// Trace: src/VX_cache_bypass.sv:28:5
					localparam MEM_TAG_ID_WIDTH = 6;
					// Trace: src/VX_cache_bypass.sv:29:5
					localparam MEM_TAG_NC1_WIDTH = 7;
					// Trace: src/VX_cache_bypass.sv:30:5
					localparam MEM_TAG_NC2_WIDTH = 7;
					// Trace: src/VX_cache_bypass.sv:31:5
					localparam MEM_TAG_OUT_WIDTH = (CACHE_ENABLE ? MEM_TAG_NC2_WIDTH : MEM_TAG_NC2_WIDTH);
					// Trace: src/VX_cache_bypass.sv:32:5
					// expanded interface instance: core_bus_nc_switch_if
					localparam _param_95306_DATA_SIZE = WORD_SIZE;
					localparam _param_95306_TAG_WIDTH = CORE_TAG_WIDTH;
					genvar _arr_95306;
					for (_arr_95306 = 0; _arr_95306 <= (((CACHE_ENABLE ? 2 : 1) * NUM_REQS) - 1); _arr_95306 = _arr_95306 + 1) begin : core_bus_nc_switch_if
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_95306_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_95306_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:7:15
						localparam UUID_WIDTH = 1;
						// Trace: src/VX_mem_bus_if.sv:9:5
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:13:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:21:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:30:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:31:5
						// Trace: src/VX_mem_bus_if.sv:39:5
					end
					// Trace: src/VX_cache_bypass.sv:36:5
					wire [0:0] core_req_nc_sel;
					// Trace: src/VX_cache_bypass.sv:37:5
					genvar _gv_i_179;
					for (_gv_i_179 = 0; _gv_i_179 < NUM_REQS; _gv_i_179 = _gv_i_179 + 1) begin : g_core_req_is_nc
						localparam i = _gv_i_179;
						if (CACHE_ENABLE) begin : g_cache
							// Trace: src/VX_cache_bypass.sv:39:13
							assign core_req_nc_sel[i] = ~Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_in_if].req_data[8];
						end
						else begin : g_no_cache
							// Trace: src/VX_cache_bypass.sv:41:13
							assign core_req_nc_sel[i] = 1'b0;
						end
					end
					// Trace: src/VX_cache_bypass.sv:44:5
					// expanded module instance: core_bus_nc_switch
					localparam _bbase_69FDB_bus_in_if = 0;
					localparam _bbase_69FDB_bus_out_if = 0;
					localparam _param_69FDB_NUM_INPUTS = NUM_REQS;
					localparam _param_69FDB_NUM_OUTPUTS = (CACHE_ENABLE ? 2 : 1) * NUM_REQS;
					localparam _param_69FDB_DATA_SIZE = WORD_SIZE;
					localparam _param_69FDB_TAG_WIDTH = CORE_TAG_WIDTH;
					localparam _param_69FDB_ARBITER = "R";
					localparam _param_69FDB_REQ_OUT_BUF = 0;
					localparam _param_69FDB_RSP_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
					if (1) begin : core_bus_nc_switch
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_switch.sv:2:15
						localparam NUM_INPUTS = _param_69FDB_NUM_INPUTS;
						// Trace: src/VX_mem_switch.sv:3:15
						localparam NUM_OUTPUTS = _param_69FDB_NUM_OUTPUTS;
						// Trace: src/VX_mem_switch.sv:4:15
						localparam DATA_SIZE = _param_69FDB_DATA_SIZE;
						// Trace: src/VX_mem_switch.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_switch.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_switch.sv:7:15
						localparam TAG_WIDTH = _param_69FDB_TAG_WIDTH;
						// Trace: src/VX_mem_switch.sv:8:15
						localparam REQ_OUT_BUF = _param_69FDB_REQ_OUT_BUF;
						// Trace: src/VX_mem_switch.sv:9:15
						localparam RSP_OUT_BUF = _param_69FDB_RSP_OUT_BUF;
						// Trace: src/VX_mem_switch.sv:10:16
						localparam ARBITER = _param_69FDB_ARBITER;
						// Trace: src/VX_mem_switch.sv:11:15
						localparam NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
						// Trace: src/VX_mem_switch.sv:12:15
						localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
						// Trace: src/VX_mem_switch.sv:13:15
						localparam LOG_NUM_REQS = $clog2(NUM_REQS);
						// Trace: src/VX_mem_switch.sv:15:5
						wire clk;
						// Trace: src/VX_mem_switch.sv:16:5
						wire reset;
						// Trace: src/VX_mem_switch.sv:17:5
						wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] bus_sel;
						// Trace: src/VX_mem_switch.sv:18:5
						localparam _mbase_bus_in_if = 0;
						// Trace: src/VX_mem_switch.sv:19:5
						localparam _mbase_bus_out_if = 0;
						// Trace: src/VX_mem_switch.sv:21:5
						localparam DATA_WIDTH = 512;
						// Trace: src/VX_mem_switch.sv:22:5
						localparam REQ_DATAW = 613;
						// Trace: src/VX_mem_switch.sv:23:5
						localparam RSP_DATAW = 519;
						// Trace: src/VX_mem_switch.sv:24:5
						wire [0:0] req_valid_in;
						// Trace: src/VX_mem_switch.sv:25:5
						wire [612:0] req_data_in;
						// Trace: src/VX_mem_switch.sv:26:5
						wire [0:0] req_ready_in;
						// Trace: src/VX_mem_switch.sv:27:5
						wire [NUM_OUTPUTS - 1:0] req_valid_out;
						// Trace: src/VX_mem_switch.sv:28:5
						wire [(NUM_OUTPUTS * 613) - 1:0] req_data_out;
						// Trace: src/VX_mem_switch.sv:29:5
						wire [NUM_OUTPUTS - 1:0] req_ready_out;
						// Trace: src/VX_mem_switch.sv:30:5
						genvar _gv_i_154;
						for (_gv_i_154 = 0; _gv_i_154 < NUM_INPUTS; _gv_i_154 = _gv_i_154 + 1) begin : g_req_data_in
							localparam i = _gv_i_154;
							// Trace: src/VX_mem_switch.sv:31:9
							assign req_valid_in[i] = Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].req_valid;
							// Trace: src/VX_mem_switch.sv:32:9
							assign req_data_in[i * 613+:613] = Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].req_data;
							// Trace: src/VX_mem_switch.sv:33:9
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
						end
						// Trace: src/VX_mem_switch.sv:35:5
						VX_stream_switch #(
							.NUM_INPUTS(NUM_INPUTS),
							.NUM_OUTPUTS(NUM_OUTPUTS),
							.DATAW(REQ_DATAW),
							.OUT_BUF(REQ_OUT_BUF)
						) req_switch(
							.clk(clk),
							.reset(reset),
							.sel_in(bus_sel),
							.valid_in(req_valid_in),
							.data_in(req_data_in),
							.ready_in(req_ready_in),
							.valid_out(req_valid_out),
							.data_out(req_data_out),
							.ready_out(req_ready_out)
						);
						// Trace: src/VX_mem_switch.sv:51:5
						genvar _gv_i_155;
						for (_gv_i_155 = 0; _gv_i_155 < NUM_OUTPUTS; _gv_i_155 = _gv_i_155 + 1) begin : g_req_data_out
							localparam i = _gv_i_155;
							// Trace: src/VX_mem_switch.sv:52:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
							// Trace: src/VX_mem_switch.sv:53:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_data = req_data_out[i * 613+:613];
							// Trace: src/VX_mem_switch.sv:54:9
							assign req_ready_out[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_ready;
						end
						// Trace: src/VX_mem_switch.sv:56:5
						wire [NUM_OUTPUTS - 1:0] rsp_valid_in;
						// Trace: src/VX_mem_switch.sv:57:5
						wire [(NUM_OUTPUTS * 519) - 1:0] rsp_data_in;
						// Trace: src/VX_mem_switch.sv:58:5
						wire [NUM_OUTPUTS - 1:0] rsp_ready_in;
						// Trace: src/VX_mem_switch.sv:59:5
						wire [0:0] rsp_valid_out;
						// Trace: src/VX_mem_switch.sv:60:5
						wire [518:0] rsp_data_out;
						// Trace: src/VX_mem_switch.sv:61:5
						wire [0:0] rsp_ready_out;
						// Trace: src/VX_mem_switch.sv:62:5
						genvar _gv_i_156;
						for (_gv_i_156 = 0; _gv_i_156 < NUM_OUTPUTS; _gv_i_156 = _gv_i_156 + 1) begin : g_rsp_data_in
							localparam i = _gv_i_156;
							// Trace: src/VX_mem_switch.sv:63:9
							assign rsp_valid_in[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_valid;
							// Trace: src/VX_mem_switch.sv:64:9
							assign rsp_data_in[i * 519+:519] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_data;
							// Trace: src/VX_mem_switch.sv:65:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
						end
						// Trace: src/VX_mem_switch.sv:67:5
						VX_stream_arb #(
							.NUM_INPUTS(NUM_OUTPUTS),
							.NUM_OUTPUTS(NUM_INPUTS),
							.DATAW(RSP_DATAW),
							.ARBITER(ARBITER),
							.OUT_BUF(RSP_OUT_BUF)
						) rsp_arb(
							.clk(clk),
							.reset(reset),
							.valid_in(rsp_valid_in),
							.data_in(rsp_data_in),
							.ready_in(rsp_ready_in),
							.valid_out(rsp_valid_out),
							.data_out(rsp_data_out),
							.ready_out(rsp_ready_out),
							.sel_out()
						);
						// Trace: src/VX_mem_switch.sv:84:5
						genvar _gv_i_157;
						for (_gv_i_157 = 0; _gv_i_157 < NUM_INPUTS; _gv_i_157 = _gv_i_157 + 1) begin : g_rsp_data_out
							localparam i = _gv_i_157;
							// Trace: src/VX_mem_switch.sv:85:9
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
							// Trace: src/VX_mem_switch.sv:86:9
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
							// Trace: src/VX_mem_switch.sv:87:9
							assign rsp_ready_out[i] = Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].rsp_ready;
						end
					end
					assign core_bus_nc_switch.clk = clk;
					assign core_bus_nc_switch.reset = reset;
					assign core_bus_nc_switch.bus_sel = core_req_nc_sel;
					// Trace: src/VX_cache_bypass.sv:59:5
					// expanded interface instance: core_bus_in_nc_if
					localparam _param_C0263_DATA_SIZE = WORD_SIZE;
					localparam _param_C0263_TAG_WIDTH = CORE_TAG_WIDTH;
					genvar _arr_C0263;
					for (_arr_C0263 = 0; _arr_C0263 <= 0; _arr_C0263 = _arr_C0263 + 1) begin : core_bus_in_nc_if
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_C0263_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_C0263_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:7:15
						localparam UUID_WIDTH = 1;
						// Trace: src/VX_mem_bus_if.sv:9:5
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:13:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:21:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:30:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:31:5
						// Trace: src/VX_mem_bus_if.sv:39:5
					end
					// Trace: src/VX_cache_bypass.sv:63:5
					genvar _gv_i_180;
					for (_gv_i_180 = 0; _gv_i_180 < NUM_REQS; _gv_i_180 = _gv_i_180 + 1) begin : g_core_bus_nc_switch_if
						localparam i = _gv_i_180;
						// Trace: src/VX_cache_bypass.sv:64:9
						assign core_bus_in_nc_if[i].req_valid = core_bus_nc_switch_if[0 + i].req_valid;
						// Trace: src/VX_cache_bypass.sv:65:9
						assign core_bus_in_nc_if[i].req_data = core_bus_nc_switch_if[0 + i].req_data;
						// Trace: src/VX_cache_bypass.sv:66:9
						assign core_bus_nc_switch_if[0 + i].req_ready = core_bus_in_nc_if[i].req_ready;
						// Trace: src/VX_cache_bypass.sv:67:9
						assign core_bus_nc_switch_if[0 + i].rsp_valid = core_bus_in_nc_if[i].rsp_valid;
						// Trace: src/VX_cache_bypass.sv:68:9
						assign core_bus_nc_switch_if[0 + i].rsp_data = core_bus_in_nc_if[i].rsp_data;
						// Trace: src/VX_cache_bypass.sv:69:9
						assign core_bus_in_nc_if[i].rsp_ready = core_bus_nc_switch_if[0 + i].rsp_ready;
						if (CACHE_ENABLE) begin : g_cache
							// Trace: src/VX_cache_bypass.sv:71:13
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = core_bus_nc_switch_if[1 + i].req_valid;
							// Trace: src/VX_cache_bypass.sv:72:13
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = core_bus_nc_switch_if[1 + i].req_data;
							// Trace: src/VX_cache_bypass.sv:73:13
							assign core_bus_nc_switch_if[1 + i].req_ready = Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_ready;
							// Trace: src/VX_cache_bypass.sv:74:13
							assign core_bus_nc_switch_if[1 + i].rsp_valid = Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_valid;
							// Trace: src/VX_cache_bypass.sv:75:13
							assign core_bus_nc_switch_if[1 + i].rsp_data = Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_data;
							// Trace: src/VX_cache_bypass.sv:76:13
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = core_bus_nc_switch_if[1 + i].rsp_ready;
						end
						else begin : g_no_cache
							// Trace: src/VX_cache_bypass.sv:78:5
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = 0;
							// Trace: src/VX_cache_bypass.sv:79:5
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = 1'sb0;
							// Trace: src/VX_cache_bypass.sv:80:5
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = 0;
						end
					end
					// Trace: src/VX_cache_bypass.sv:83:5
					// expanded interface instance: core_bus_nc_arb_if
					localparam _param_D50AC_DATA_SIZE = WORD_SIZE;
					localparam _param_D50AC_TAG_WIDTH = MEM_TAG_NC1_WIDTH;
					genvar _arr_D50AC;
					for (_arr_D50AC = 0; _arr_D50AC <= 0; _arr_D50AC = _arr_D50AC + 1) begin : core_bus_nc_arb_if
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_D50AC_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_D50AC_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:7:15
						localparam UUID_WIDTH = 1;
						// Trace: src/VX_mem_bus_if.sv:9:5
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:13:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:21:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:30:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:31:5
						// Trace: src/VX_mem_bus_if.sv:39:5
					end
					// Trace: src/VX_cache_bypass.sv:87:5
					// expanded module instance: core_bus_nc_arb
					localparam _bbase_1376F_bus_in_if = 0;
					localparam _bbase_1376F_bus_out_if = 0;
					localparam _param_1376F_NUM_INPUTS = NUM_REQS;
					localparam _param_1376F_NUM_OUTPUTS = MEM_PORTS;
					localparam _param_1376F_DATA_SIZE = WORD_SIZE;
					localparam _param_1376F_TAG_WIDTH = CORE_TAG_WIDTH;
					localparam _param_1376F_TAG_SEL_IDX = TAG_SEL_IDX;
					localparam _param_1376F_ARBITER = (CACHE_ENABLE ? "P" : "R");
					localparam _param_1376F_REQ_OUT_BUF = 0;
					localparam _param_1376F_RSP_OUT_BUF = 0;
					if (1) begin : core_bus_nc_arb
						// Trace: src/VX_mem_arb.sv:2:15
						localparam NUM_INPUTS = _param_1376F_NUM_INPUTS;
						// Trace: src/VX_mem_arb.sv:3:15
						localparam NUM_OUTPUTS = _param_1376F_NUM_OUTPUTS;
						// Trace: src/VX_mem_arb.sv:4:15
						localparam DATA_SIZE = _param_1376F_DATA_SIZE;
						// Trace: src/VX_mem_arb.sv:5:15
						localparam TAG_WIDTH = _param_1376F_TAG_WIDTH;
						// Trace: src/VX_mem_arb.sv:6:15
						localparam TAG_SEL_IDX = _param_1376F_TAG_SEL_IDX;
						// Trace: src/VX_mem_arb.sv:7:15
						localparam REQ_OUT_BUF = _param_1376F_REQ_OUT_BUF;
						// Trace: src/VX_mem_arb.sv:8:15
						localparam RSP_OUT_BUF = _param_1376F_RSP_OUT_BUF;
						// Trace: src/VX_mem_arb.sv:9:16
						localparam ARBITER = _param_1376F_ARBITER;
						// Trace: src/VX_mem_arb.sv:10:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_arb.sv:11:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_arb.sv:12:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_arb.sv:14:5
						wire clk;
						// Trace: src/VX_mem_arb.sv:15:5
						wire reset;
						// Trace: src/VX_mem_arb.sv:16:5
						localparam _mbase_bus_in_if = 0;
						// Trace: src/VX_mem_arb.sv:17:5
						localparam _mbase_bus_out_if = 0;
						// Trace: src/VX_mem_arb.sv:19:5
						localparam DATA_WIDTH = 512;
						// Trace: src/VX_mem_arb.sv:20:5
						localparam LOG_NUM_REQS = 0;
						// Trace: src/VX_mem_arb.sv:21:5
						localparam REQ_DATAW = 613;
						// Trace: src/VX_mem_arb.sv:22:5
						localparam RSP_DATAW = 519;
						// Trace: src/VX_mem_arb.sv:24:5
						wire [0:0] req_valid_in;
						// Trace: src/VX_mem_arb.sv:25:5
						wire [612:0] req_data_in;
						// Trace: src/VX_mem_arb.sv:26:5
						wire [0:0] req_ready_in;
						// Trace: src/VX_mem_arb.sv:27:5
						wire [0:0] req_valid_out;
						// Trace: src/VX_mem_arb.sv:28:5
						wire [612:0] req_data_out;
						// Trace: src/VX_mem_arb.sv:29:5
						wire [0:0] req_sel_out;
						// Trace: src/VX_mem_arb.sv:30:5
						wire [0:0] req_ready_out;
						// Trace: src/VX_mem_arb.sv:31:5
						genvar _gv_i_80;
						for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
							localparam i = _gv_i_80;
							// Trace: src/VX_mem_arb.sv:32:9
							assign req_valid_in[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_valid;
							// Trace: src/VX_mem_arb.sv:33:9
							assign req_data_in[i * 613+:613] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_data;
							// Trace: src/VX_mem_arb.sv:34:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
						end
						// Trace: src/VX_mem_arb.sv:36:5
						VX_stream_arb #(
							.NUM_INPUTS(NUM_INPUTS),
							.NUM_OUTPUTS(NUM_OUTPUTS),
							.DATAW(REQ_DATAW),
							.ARBITER(ARBITER),
							.OUT_BUF(REQ_OUT_BUF)
						) req_arb(
							.clk(clk),
							.reset(reset),
							.valid_in(req_valid_in),
							.ready_in(req_ready_in),
							.data_in(req_data_in),
							.data_out(req_data_out),
							.sel_out(req_sel_out),
							.valid_out(req_valid_out),
							.ready_out(req_ready_out)
						);
						// Trace: src/VX_mem_arb.sv:53:5
						genvar _gv_i_81;
						for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
							localparam i = _gv_i_81;
							// Trace: src/VX_mem_arb.sv:54:9
							wire [6:0] req_tag_out;
							// Trace: src/VX_mem_arb.sv:55:9
							VX_bits_insert #(
								.N(TAG_WIDTH),
								.S(LOG_NUM_REQS),
								.POS(TAG_SEL_IDX)
							) bits_insert(
								.data_in(req_tag_out),
								.ins_in(req_sel_out[i+:1]),
								.data_out(Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[6-:7])
							);
							// Trace: src/VX_mem_arb.sv:64:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
							// Trace: src/VX_mem_arb.sv:65:9
							assign {Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[612], Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[611-:26], Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[585-:512], Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[73-:64], Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[9-:3], req_tag_out} = req_data_out[i * 613+:613];
							// Trace: src/VX_mem_arb.sv:73:9
							assign req_ready_out[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_ready;
						end
						// Trace: src/VX_mem_arb.sv:75:5
						wire [0:0] rsp_valid_out;
						// Trace: src/VX_mem_arb.sv:76:5
						wire [518:0] rsp_data_out;
						// Trace: src/VX_mem_arb.sv:77:5
						wire [0:0] rsp_ready_out;
						// Trace: src/VX_mem_arb.sv:78:5
						wire [0:0] rsp_valid_in;
						// Trace: src/VX_mem_arb.sv:79:5
						wire [518:0] rsp_data_in;
						// Trace: src/VX_mem_arb.sv:80:5
						wire [0:0] rsp_ready_in;
						// Trace: src/VX_mem_arb.sv:81:5
						if (1) begin : g_passthru
							genvar _gv_i_83;
							for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
								localparam i = _gv_i_83;
								// Trace: src/VX_mem_arb.sv:116:13
								assign rsp_valid_in[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_valid;
								// Trace: src/VX_mem_arb.sv:117:13
								assign rsp_data_in[i * 519+:519] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_data;
								// Trace: src/VX_mem_arb.sv:118:13
								assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
							end
							// Trace: src/VX_mem_arb.sv:120:9
							VX_stream_arb #(
								.NUM_INPUTS(NUM_OUTPUTS),
								.NUM_OUTPUTS(NUM_INPUTS),
								.DATAW(RSP_DATAW),
								.ARBITER(ARBITER),
								.OUT_BUF(RSP_OUT_BUF)
							) req_arb(
								.clk(clk),
								.reset(reset),
								.valid_in(rsp_valid_in),
								.ready_in(rsp_ready_in),
								.data_in(rsp_data_in),
								.data_out(rsp_data_out),
								.valid_out(rsp_valid_out),
								.ready_out(rsp_ready_out),
								.sel_out()
							);
						end
						// Trace: src/VX_mem_arb.sv:138:5
						genvar _gv_i_84;
						for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
							localparam i = _gv_i_84;
							// Trace: src/VX_mem_arb.sv:139:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
							// Trace: src/VX_mem_arb.sv:140:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
							// Trace: src/VX_mem_arb.sv:141:9
							assign rsp_ready_out[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_ready;
						end
					end
					assign core_bus_nc_arb.clk = clk;
					assign core_bus_nc_arb.reset = reset;
					// Trace: src/VX_cache_bypass.sv:102:5
					// expanded interface instance: mem_bus_out_nc_if
					localparam _param_0061C_DATA_SIZE = LINE_SIZE;
					localparam _param_0061C_TAG_WIDTH = MEM_TAG_NC2_WIDTH;
					genvar _arr_0061C;
					for (_arr_0061C = 0; _arr_0061C <= 0; _arr_0061C = _arr_0061C + 1) begin : mem_bus_out_nc_if
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_0061C_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_0061C_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:7:15
						localparam UUID_WIDTH = 1;
						// Trace: src/VX_mem_bus_if.sv:9:5
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:13:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:21:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:30:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:31:5
						// Trace: src/VX_mem_bus_if.sv:39:5
					end
					// Trace: src/VX_cache_bypass.sv:106:5
					genvar _gv_i_181;
					for (_gv_i_181 = 0; _gv_i_181 < MEM_PORTS; _gv_i_181 = _gv_i_181 + 1) begin : g_mem_bus_out_nc
						localparam i = _gv_i_181;
						// Trace: src/VX_cache_bypass.sv:107:9
						wire core_req_nc_arb_rw;
						// Trace: src/VX_cache_bypass.sv:108:9
						wire [63:0] core_req_nc_arb_byteen;
						// Trace: src/VX_cache_bypass.sv:109:9
						wire [25:0] core_req_nc_arb_addr;
						// Trace: src/VX_cache_bypass.sv:110:9
						wire [2:0] core_req_nc_arb_flags;
						// Trace: src/VX_cache_bypass.sv:111:9
						wire [511:0] core_req_nc_arb_data;
						// Trace: src/VX_cache_bypass.sv:112:9
						wire [6:0] core_req_nc_arb_tag;
						// Trace: src/VX_cache_bypass.sv:113:9
						assign {core_req_nc_arb_rw, core_req_nc_arb_addr, core_req_nc_arb_data, core_req_nc_arb_byteen, core_req_nc_arb_flags, core_req_nc_arb_tag} = core_bus_nc_arb_if[i].req_data;
						// Trace: src/VX_cache_bypass.sv:121:9
						wire [25:0] core_req_nc_arb_addr_w;
						// Trace: src/VX_cache_bypass.sv:122:9
						wire [63:0] core_req_nc_arb_byteen_w;
						// Trace: src/VX_cache_bypass.sv:123:9
						wire [511:0] core_req_nc_arb_data_w;
						// Trace: src/VX_cache_bypass.sv:124:9
						wire [511:0] core_rsp_nc_arb_data_w;
						// Trace: src/VX_cache_bypass.sv:125:9
						wire [6:0] core_req_nc_arb_tag_w;
						// Trace: src/VX_cache_bypass.sv:126:9
						wire [6:0] core_rsp_nc_arb_tag_w;
						if (1) begin : g_single_word_line
							// Trace: src/VX_cache_bypass.sv:157:13
							assign core_req_nc_arb_addr_w = core_req_nc_arb_addr;
							// Trace: src/VX_cache_bypass.sv:158:13
							assign core_req_nc_arb_byteen_w = core_req_nc_arb_byteen;
							// Trace: src/VX_cache_bypass.sv:159:13
							assign core_req_nc_arb_data_w = core_req_nc_arb_data;
							// Trace: src/VX_cache_bypass.sv:160:13
							assign core_req_nc_arb_tag_w = core_req_nc_arb_tag;
							// Trace: src/VX_cache_bypass.sv:161:13
							assign core_rsp_nc_arb_data_w = mem_bus_out_nc_if[i].rsp_data[518-:512];
							// Trace: src/VX_cache_bypass.sv:162:13
							assign core_rsp_nc_arb_tag_w = sv2v_cast_7(mem_bus_out_nc_if[i].rsp_data[6-:7]);
						end
						// Trace: src/VX_cache_bypass.sv:164:9
						assign mem_bus_out_nc_if[i].req_valid = core_bus_nc_arb_if[i].req_valid;
						// Trace: src/VX_cache_bypass.sv:165:9
						assign mem_bus_out_nc_if[i].req_data = {core_req_nc_arb_rw, core_req_nc_arb_addr_w, core_req_nc_arb_data_w, core_req_nc_arb_byteen_w, core_req_nc_arb_flags, core_req_nc_arb_tag_w};
						// Trace: src/VX_cache_bypass.sv:173:9
						assign core_bus_nc_arb_if[i].req_ready = mem_bus_out_nc_if[i].req_ready;
						// Trace: src/VX_cache_bypass.sv:174:9
						assign core_bus_nc_arb_if[i].rsp_valid = mem_bus_out_nc_if[i].rsp_valid;
						// Trace: src/VX_cache_bypass.sv:175:9
						assign core_bus_nc_arb_if[i].rsp_data = {core_rsp_nc_arb_data_w, core_rsp_nc_arb_tag_w};
						// Trace: src/VX_cache_bypass.sv:179:9
						assign mem_bus_out_nc_if[i].rsp_ready = core_bus_nc_arb_if[i].rsp_ready;
					end
					// Trace: src/VX_cache_bypass.sv:181:5
					// expanded interface instance: mem_bus_out_src_if
					localparam _param_913F6_DATA_SIZE = LINE_SIZE;
					localparam _param_913F6_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
					genvar _arr_913F6;
					for (_arr_913F6 = 0; _arr_913F6 <= (((CACHE_ENABLE ? 2 : 1) * MEM_PORTS) - 1); _arr_913F6 = _arr_913F6 + 1) begin : mem_bus_out_src_if
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_913F6_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_913F6_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:7:15
						localparam UUID_WIDTH = 1;
						// Trace: src/VX_mem_bus_if.sv:9:5
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:13:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:21:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire [(606 + (_param_913F6_TAG_WIDTH + 0)) - 1:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire [(512 + (_param_913F6_TAG_WIDTH + 0)) - 1:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:30:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:31:5
						// Trace: src/VX_mem_bus_if.sv:39:5
					end
					// Trace: src/VX_cache_bypass.sv:185:5
					genvar _gv_i_182;
					for (_gv_i_182 = 0; _gv_i_182 < MEM_PORTS; _gv_i_182 = _gv_i_182 + 1) begin : g_mem_bus_out_src
						localparam i = _gv_i_182;
						// Trace: src/VX_cache_bypass.sv:186:5
						assign mem_bus_out_src_if[0 + i].req_valid = mem_bus_out_nc_if[i].req_valid;
						// Trace: src/VX_cache_bypass.sv:187:5
						assign mem_bus_out_src_if[0 + i].req_data[539 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))] = mem_bus_out_nc_if[i].req_data[612];
						// Trace: src/VX_cache_bypass.sv:188:5
						assign mem_bus_out_src_if[0 + i].req_data[538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))-:((602 + (_param_913F6_TAG_WIDTH + 2)) >= (579 + (_param_913F6_TAG_WIDTH + 0)) ? ((538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) - (512 + (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0))))) + 1 : ((512 + (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0)))) - (538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)))) + 1)] = mem_bus_out_nc_if[i].req_data[611-:26];
						// Trace: src/VX_cache_bypass.sv:189:5
						assign mem_bus_out_src_if[0 + i].req_data[512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))-:((576 + (_param_913F6_TAG_WIDTH + 2)) >= (67 + (_param_913F6_TAG_WIDTH + 0)) ? ((512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) - (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0)))) + 1 : ((_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0))) - (512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)))) + 1)] = mem_bus_out_nc_if[i].req_data[585-:512];
						// Trace: src/VX_cache_bypass.sv:190:5
						assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)-:((_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)) >= (3 + (_param_913F6_TAG_WIDTH + 0)) ? ((_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)) - (3 + (_param_913F6_TAG_WIDTH + 0))) + 1 : ((3 + (_param_913F6_TAG_WIDTH + 0)) - (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) + 1)] = mem_bus_out_nc_if[i].req_data[73-:64];
						// Trace: src/VX_cache_bypass.sv:191:5
						assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_TAG_WIDTH + 2-:((_param_913F6_TAG_WIDTH + 2) >= (_param_913F6_TAG_WIDTH + 0) ? ((_param_913F6_TAG_WIDTH + 2) - (_param_913F6_TAG_WIDTH + 0)) + 1 : ((_param_913F6_TAG_WIDTH + 0) - (_param_913F6_TAG_WIDTH + 2)) + 1)] = mem_bus_out_nc_if[i].req_data[9-:3];
						if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk1
							if (1) begin : genblk1
								if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
									// Trace: src/VX_cache_bypass.sv:196:17
									assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = {mem_bus_out_nc_if[i].req_data[6-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_NC2_WIDTH {1'b0}}, mem_bus_out_nc_if[i].req_data[5-:6]};
								end
								else begin : genblk1
									// Trace: src/VX_cache_bypass.sv:198:17
									assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = {mem_bus_out_nc_if[i].req_data[6-:1], mem_bus_out_nc_if[i].req_data[6 - (1 + (6 - (MEM_TAG_OUT_WIDTH - UUID_WIDTH))):0]};
								end
							end
						end
						else begin : genblk1
							// Trace: src/VX_cache_bypass.sv:208:9
							assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = mem_bus_out_nc_if[i].req_data[6-:7];
						end
						// Trace: src/VX_cache_bypass.sv:211:5
						assign mem_bus_out_nc_if[i].req_ready = mem_bus_out_src_if[0 + i].req_ready;
						// Trace: src/VX_cache_bypass.sv:212:5
						assign mem_bus_out_nc_if[i].rsp_valid = mem_bus_out_src_if[0 + i].rsp_valid;
						// Trace: src/VX_cache_bypass.sv:213:5
						assign mem_bus_out_nc_if[i].rsp_data[518-:512] = mem_bus_out_src_if[0 + i].rsp_data[_param_913F6_TAG_WIDTH + 511-:((_param_913F6_TAG_WIDTH + 511) >= (_param_913F6_TAG_WIDTH + 0) ? ((_param_913F6_TAG_WIDTH + 511) - (_param_913F6_TAG_WIDTH + 0)) + 1 : ((_param_913F6_TAG_WIDTH + 0) - (_param_913F6_TAG_WIDTH + 511)) + 1)];
						if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk2
							if (1) begin : genblk1
								if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
									// Trace: src/VX_cache_bypass.sv:218:17
									assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1))-:((_param_913F6_TAG_WIDTH - 1) >= (_param_913F6_TAG_WIDTH - 1) ? ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1 : ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1)], mem_bus_out_src_if[0 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 2) - (_param_913F6_TAG_WIDTH - 7))):(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 2) - (_param_913F6_TAG_WIDTH - 2)))]};
								end
								else begin : genblk1
									// Trace: src/VX_cache_bypass.sv:220:17
									assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1))-:((_param_913F6_TAG_WIDTH - 1) >= (_param_913F6_TAG_WIDTH - 1) ? ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1 : ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1)], {MEM_TAG_NC2_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[0 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 2))-:_param_913F6_TAG_WIDTH - 1]};
								end
							end
						end
						else begin : genblk2
							// Trace: src/VX_cache_bypass.sv:230:9
							assign mem_bus_out_nc_if[i].rsp_data[6-:7] = mem_bus_out_src_if[0 + i].rsp_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0];
						end
						// Trace: src/VX_cache_bypass.sv:233:5
						assign mem_bus_out_src_if[0 + i].rsp_ready = mem_bus_out_nc_if[i].rsp_ready;
						if (CACHE_ENABLE) begin : g_cache
							// Trace: src/VX_cache_bypass.sv:235:5
							assign mem_bus_out_src_if[1 + i].req_valid = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_valid;
							// Trace: src/VX_cache_bypass.sv:236:5
							assign mem_bus_out_src_if[1 + i].req_data[539 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[610];
							// Trace: src/VX_cache_bypass.sv:237:5
							assign mem_bus_out_src_if[1 + i].req_data[538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))-:((602 + (_param_913F6_TAG_WIDTH + 2)) >= (579 + (_param_913F6_TAG_WIDTH + 0)) ? ((538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) - (512 + (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0))))) + 1 : ((512 + (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0)))) - (538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)))) + 1)] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[609-:26];
							// Trace: src/VX_cache_bypass.sv:238:5
							assign mem_bus_out_src_if[1 + i].req_data[512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))-:((576 + (_param_913F6_TAG_WIDTH + 2)) >= (67 + (_param_913F6_TAG_WIDTH + 0)) ? ((512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) - (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0)))) + 1 : ((_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0))) - (512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)))) + 1)] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[583-:512];
							// Trace: src/VX_cache_bypass.sv:239:5
							assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)-:((_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)) >= (3 + (_param_913F6_TAG_WIDTH + 0)) ? ((_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)) - (3 + (_param_913F6_TAG_WIDTH + 0))) + 1 : ((3 + (_param_913F6_TAG_WIDTH + 0)) - (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) + 1)] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[71-:64];
							// Trace: src/VX_cache_bypass.sv:240:5
							assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_TAG_WIDTH + 2-:((_param_913F6_TAG_WIDTH + 2) >= (_param_913F6_TAG_WIDTH + 0) ? ((_param_913F6_TAG_WIDTH + 2) - (_param_913F6_TAG_WIDTH + 0)) + 1 : ((_param_913F6_TAG_WIDTH + 0) - (_param_913F6_TAG_WIDTH + 2)) + 1)] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[7-:3];
							if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk1
								if (1) begin : genblk1
									if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
										// Trace: src/VX_cache_bypass.sv:245:17
										assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = {Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_IN_WIDTH {1'b0}}, Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[3-:4]};
									end
									else begin : genblk1
										// Trace: src/VX_cache_bypass.sv:247:17
										assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = {Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4 - (1 + (4 - (MEM_TAG_OUT_WIDTH - UUID_WIDTH))):0]};
									end
								end
							end
							else begin : genblk1
								// Trace: src/VX_cache_bypass.sv:257:9
								assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:5];
							end
							// Trace: src/VX_cache_bypass.sv:260:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = mem_bus_out_src_if[1 + i].req_ready;
							// Trace: src/VX_cache_bypass.sv:261:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = mem_bus_out_src_if[1 + i].rsp_valid;
							// Trace: src/VX_cache_bypass.sv:262:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[516-:512] = mem_bus_out_src_if[1 + i].rsp_data[_param_913F6_TAG_WIDTH + 511-:((_param_913F6_TAG_WIDTH + 511) >= (_param_913F6_TAG_WIDTH + 0) ? ((_param_913F6_TAG_WIDTH + 511) - (_param_913F6_TAG_WIDTH + 0)) + 1 : ((_param_913F6_TAG_WIDTH + 0) - (_param_913F6_TAG_WIDTH + 511)) + 1)];
							if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk2
								if (1) begin : genblk1
									if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
										// Trace: src/VX_cache_bypass.sv:267:17
										assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1))-:((_param_913F6_TAG_WIDTH - 1) >= (_param_913F6_TAG_WIDTH - 1) ? ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1 : ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1)], mem_bus_out_src_if[1 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 2) - (_param_913F6_TAG_WIDTH - 5))):(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 2) - (_param_913F6_TAG_WIDTH - 2)))]};
									end
									else begin : genblk1
										// Trace: src/VX_cache_bypass.sv:269:17
										assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1))-:((_param_913F6_TAG_WIDTH - 1) >= (_param_913F6_TAG_WIDTH - 1) ? ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1 : ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1)], {MEM_TAG_IN_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[1 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 2))-:_param_913F6_TAG_WIDTH - 1]};
									end
								end
							end
							else begin : genblk2
								// Trace: src/VX_cache_bypass.sv:279:9
								assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = mem_bus_out_src_if[1 + i].rsp_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0];
							end
							// Trace: src/VX_cache_bypass.sv:282:5
							assign mem_bus_out_src_if[1 + i].rsp_ready = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_ready;
						end
						else begin : g_no_cache
							// Trace: src/VX_cache_bypass.sv:284:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = 0;
							// Trace: src/VX_cache_bypass.sv:285:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = 0;
							// Trace: src/VX_cache_bypass.sv:286:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data = 1'sb0;
						end
					end
					// Trace: src/VX_cache_bypass.sv:289:5
					// expanded module instance: mem_bus_out_arb
					localparam _bbase_B06D0_bus_in_if = 0;
					localparam _bbase_B06D0_bus_out_if = 0;
					localparam _param_B06D0_NUM_INPUTS = (CACHE_ENABLE ? 2 : 1) * MEM_PORTS;
					localparam _param_B06D0_NUM_OUTPUTS = MEM_PORTS;
					localparam _param_B06D0_DATA_SIZE = LINE_SIZE;
					localparam _param_B06D0_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
					localparam _param_B06D0_ARBITER = "R";
					localparam _param_B06D0_REQ_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
					localparam _param_B06D0_RSP_OUT_BUF = 0;
					if (1) begin : mem_bus_out_arb
						// Trace: src/VX_mem_arb.sv:2:15
						localparam NUM_INPUTS = _param_B06D0_NUM_INPUTS;
						// Trace: src/VX_mem_arb.sv:3:15
						localparam NUM_OUTPUTS = _param_B06D0_NUM_OUTPUTS;
						// Trace: src/VX_mem_arb.sv:4:15
						localparam DATA_SIZE = _param_B06D0_DATA_SIZE;
						// Trace: src/VX_mem_arb.sv:5:15
						localparam TAG_WIDTH = _param_B06D0_TAG_WIDTH;
						// Trace: src/VX_mem_arb.sv:6:15
						localparam TAG_SEL_IDX = 0;
						// Trace: src/VX_mem_arb.sv:7:15
						localparam REQ_OUT_BUF = _param_B06D0_REQ_OUT_BUF;
						// Trace: src/VX_mem_arb.sv:8:15
						localparam RSP_OUT_BUF = _param_B06D0_RSP_OUT_BUF;
						// Trace: src/VX_mem_arb.sv:9:16
						localparam ARBITER = _param_B06D0_ARBITER;
						// Trace: src/VX_mem_arb.sv:10:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_arb.sv:11:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_arb.sv:12:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_arb.sv:14:5
						wire clk;
						// Trace: src/VX_mem_arb.sv:15:5
						wire reset;
						// Trace: src/VX_mem_arb.sv:16:5
						localparam _mbase_bus_in_if = 0;
						// Trace: src/VX_mem_arb.sv:17:5
						localparam _mbase_bus_out_if = 0;
						// Trace: src/VX_mem_arb.sv:19:5
						localparam DATA_WIDTH = 512;
						// Trace: src/VX_mem_arb.sv:20:5
						localparam LOG_NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? $clog2((NUM_INPUTS + 0) / 1) : 0);
						// Trace: src/VX_mem_arb.sv:21:5
						localparam REQ_DATAW = 606 + TAG_WIDTH;
						// Trace: src/VX_mem_arb.sv:22:5
						localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
						// Trace: src/VX_mem_arb.sv:24:5
						wire [NUM_INPUTS - 1:0] req_valid_in;
						// Trace: src/VX_mem_arb.sv:25:5
						wire [(NUM_INPUTS * REQ_DATAW) - 1:0] req_data_in;
						// Trace: src/VX_mem_arb.sv:26:5
						wire [NUM_INPUTS - 1:0] req_ready_in;
						// Trace: src/VX_mem_arb.sv:27:5
						wire [0:0] req_valid_out;
						// Trace: src/VX_mem_arb.sv:28:5
						wire [REQ_DATAW - 1:0] req_data_out;
						// Trace: src/VX_mem_arb.sv:29:5
						wire [(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1) - 1:0] req_sel_out;
						// Trace: src/VX_mem_arb.sv:30:5
						wire [0:0] req_ready_out;
						// Trace: src/VX_mem_arb.sv:31:5
						genvar _gv_i_80;
						for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
							localparam i = _gv_i_80;
							// Trace: src/VX_mem_arb.sv:32:9
							assign req_valid_in[i] = Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_valid;
							// Trace: src/VX_mem_arb.sv:33:9
							assign req_data_in[i * REQ_DATAW+:REQ_DATAW] = Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_data;
							// Trace: src/VX_mem_arb.sv:34:9
							assign Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
						end
						// Trace: src/VX_mem_arb.sv:36:5
						VX_stream_arb #(
							.NUM_INPUTS(NUM_INPUTS),
							.NUM_OUTPUTS(NUM_OUTPUTS),
							.DATAW(REQ_DATAW),
							.ARBITER(ARBITER),
							.OUT_BUF(REQ_OUT_BUF)
						) req_arb(
							.clk(clk),
							.reset(reset),
							.valid_in(req_valid_in),
							.ready_in(req_ready_in),
							.data_in(req_data_in),
							.data_out(req_data_out),
							.sel_out(req_sel_out),
							.valid_out(req_valid_out),
							.ready_out(req_ready_out)
						);
						// Trace: src/VX_mem_arb.sv:53:5
						genvar _gv_i_81;
						for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
							localparam i = _gv_i_81;
							// Trace: src/VX_mem_arb.sv:54:9
							wire [TAG_WIDTH - 1:0] req_tag_out;
							// Trace: src/VX_mem_arb.sv:55:9
							VX_bits_insert #(
								.N(TAG_WIDTH),
								.S(LOG_NUM_REQS),
								.POS(TAG_SEL_IDX)
							) bits_insert(
								.data_in(req_tag_out),
								.ins_in(req_sel_out[i * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)]),
								.data_out(Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[_param_4FE36_TAG_WIDTH - 1-:_param_4FE36_TAG_WIDTH + 0])
							);
							// Trace: src/VX_mem_arb.sv:64:9
							assign Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
							// Trace: src/VX_mem_arb.sv:65:9
							assign {Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[539 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))], Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))-:((602 + (_param_4FE36_TAG_WIDTH + 2)) >= (579 + (_param_4FE36_TAG_WIDTH + 0)) ? ((538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))) - (512 + (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0))))) + 1 : ((512 + (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0)))) - (538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)))) + 1)], Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[512 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))-:((576 + (_param_4FE36_TAG_WIDTH + 2)) >= (67 + (_param_4FE36_TAG_WIDTH + 0)) ? ((512 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))) - (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0)))) + 1 : ((_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0))) - (512 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)))) + 1)], Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)-:((_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)) >= (3 + (_param_4FE36_TAG_WIDTH + 0)) ? ((_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)) - (3 + (_param_4FE36_TAG_WIDTH + 0))) + 1 : ((3 + (_param_4FE36_TAG_WIDTH + 0)) - (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))) + 1)], Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[_param_4FE36_TAG_WIDTH + 2-:((_param_4FE36_TAG_WIDTH + 2) >= (_param_4FE36_TAG_WIDTH + 0) ? ((_param_4FE36_TAG_WIDTH + 2) - (_param_4FE36_TAG_WIDTH + 0)) + 1 : ((_param_4FE36_TAG_WIDTH + 0) - (_param_4FE36_TAG_WIDTH + 2)) + 1)], req_tag_out} = req_data_out[i * REQ_DATAW+:REQ_DATAW];
							// Trace: src/VX_mem_arb.sv:73:9
							assign req_ready_out[i] = Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
						end
						// Trace: src/VX_mem_arb.sv:75:5
						wire [NUM_INPUTS - 1:0] rsp_valid_out;
						// Trace: src/VX_mem_arb.sv:76:5
						wire [(NUM_INPUTS * RSP_DATAW) - 1:0] rsp_data_out;
						// Trace: src/VX_mem_arb.sv:77:5
						wire [NUM_INPUTS - 1:0] rsp_ready_out;
						// Trace: src/VX_mem_arb.sv:78:5
						wire [0:0] rsp_valid_in;
						// Trace: src/VX_mem_arb.sv:79:5
						wire [RSP_DATAW - 1:0] rsp_data_in;
						// Trace: src/VX_mem_arb.sv:80:5
						wire [0:0] rsp_ready_in;
						// Trace: src/VX_mem_arb.sv:81:5
						if (NUM_INPUTS > NUM_OUTPUTS) begin : g_rsp_enabled
							// Trace: src/VX_mem_arb.sv:82:9
							wire [LOG_NUM_REQS - 1:0] rsp_sel_in;
							genvar _gv_i_82;
							for (_gv_i_82 = 0; _gv_i_82 < NUM_OUTPUTS; _gv_i_82 = _gv_i_82 + 1) begin : g_rsp_data_in
								localparam i = _gv_i_82;
								// Trace: src/VX_mem_arb.sv:84:13
								wire [TAG_WIDTH - 1:0] rsp_tag_out;
								// Trace: src/VX_mem_arb.sv:85:13
								VX_bits_remove #(
									.N(TAG_WIDTH + LOG_NUM_REQS),
									.S(LOG_NUM_REQS),
									.POS(TAG_SEL_IDX)
								) bits_remove(
									.data_in(Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[_param_4FE36_TAG_WIDTH - 1-:_param_4FE36_TAG_WIDTH + 0]),
									.sel_out(rsp_sel_in[i * LOG_NUM_REQS+:LOG_NUM_REQS]),
									.data_out(rsp_tag_out)
								);
								// Trace: src/VX_mem_arb.sv:94:13
								assign rsp_valid_in[i] = Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
								// Trace: src/VX_mem_arb.sv:95:13
								assign rsp_data_in[i * RSP_DATAW+:RSP_DATAW] = {Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[_param_4FE36_TAG_WIDTH + 511-:((_param_4FE36_TAG_WIDTH + 511) >= (_param_4FE36_TAG_WIDTH + 0) ? ((_param_4FE36_TAG_WIDTH + 511) - (_param_4FE36_TAG_WIDTH + 0)) + 1 : ((_param_4FE36_TAG_WIDTH + 0) - (_param_4FE36_TAG_WIDTH + 511)) + 1)], rsp_tag_out};
								// Trace: src/VX_mem_arb.sv:96:13
								assign Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
							end
							// Trace: src/VX_mem_arb.sv:98:9
							VX_stream_switch #(
								.NUM_INPUTS(NUM_OUTPUTS),
								.NUM_OUTPUTS(NUM_INPUTS),
								.DATAW(RSP_DATAW),
								.OUT_BUF(RSP_OUT_BUF)
							) rsp_switch(
								.clk(clk),
								.reset(reset),
								.sel_in(rsp_sel_in),
								.valid_in(rsp_valid_in),
								.ready_in(rsp_ready_in),
								.data_in(rsp_data_in),
								.data_out(rsp_data_out),
								.valid_out(rsp_valid_out),
								.ready_out(rsp_ready_out)
							);
						end
						else begin : g_passthru
							genvar _gv_i_83;
							for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
								localparam i = _gv_i_83;
								// Trace: src/VX_mem_arb.sv:116:13
								assign rsp_valid_in[i] = Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
								// Trace: src/VX_mem_arb.sv:117:13
								assign rsp_data_in[i * RSP_DATAW+:RSP_DATAW] = Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
								// Trace: src/VX_mem_arb.sv:118:13
								assign Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
							end
							// Trace: src/VX_mem_arb.sv:120:9
							VX_stream_arb #(
								.NUM_INPUTS(NUM_OUTPUTS),
								.NUM_OUTPUTS(NUM_INPUTS),
								.DATAW(RSP_DATAW),
								.ARBITER(ARBITER),
								.OUT_BUF(RSP_OUT_BUF)
							) req_arb(
								.clk(clk),
								.reset(reset),
								.valid_in(rsp_valid_in),
								.ready_in(rsp_ready_in),
								.data_in(rsp_data_in),
								.data_out(rsp_data_out),
								.valid_out(rsp_valid_out),
								.ready_out(rsp_ready_out),
								.sel_out()
							);
						end
						// Trace: src/VX_mem_arb.sv:138:5
						genvar _gv_i_84;
						for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
							localparam i = _gv_i_84;
							// Trace: src/VX_mem_arb.sv:139:9
							assign Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
							// Trace: src/VX_mem_arb.sv:140:9
							assign Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * RSP_DATAW+:RSP_DATAW];
							// Trace: src/VX_mem_arb.sv:141:9
							assign rsp_ready_out[i] = Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_ready;
						end
					end
					assign mem_bus_out_arb.clk = clk;
					assign mem_bus_out_arb.reset = reset;
				end
				assign cache_bypass.clk = clk;
				assign cache_bypass.reset = reset;
			end
			else begin : g_no_bypass
				genvar _gv_i_167;
				for (_gv_i_167 = 0; _gv_i_167 < NUM_REQS; _gv_i_167 = _gv_i_167 + 1) begin : g_core_bus_cache_if
					localparam i = _gv_i_167;
					// Trace: src/VX_cache_wrap.sv:76:5
					assign core_bus_cache_if[i].req_valid = Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].req_valid;
					// Trace: src/VX_cache_wrap.sv:77:5
					assign core_bus_cache_if[i].req_data = Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].req_data;
					// Trace: src/VX_cache_wrap.sv:78:5
					assign Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].req_ready = core_bus_cache_if[i].req_ready;
					// Trace: src/VX_cache_wrap.sv:79:5
					assign Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].rsp_valid = core_bus_cache_if[i].rsp_valid;
					// Trace: src/VX_cache_wrap.sv:80:5
					assign Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].rsp_data = core_bus_cache_if[i].rsp_data;
					// Trace: src/VX_cache_wrap.sv:81:5
					assign core_bus_cache_if[i].rsp_ready = Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].rsp_ready;
				end
				genvar _gv_i_168;
				for (_gv_i_168 = 0; _gv_i_168 < MEM_PORTS; _gv_i_168 = _gv_i_168 + 1) begin : g_mem_bus_tmp_if
					localparam i = _gv_i_168;
					// Trace: src/VX_cache_wrap.sv:84:5
					assign mem_bus_tmp_if[i].req_valid = mem_bus_cache_if[i].req_valid;
					// Trace: src/VX_cache_wrap.sv:85:5
					assign mem_bus_tmp_if[i].req_data = mem_bus_cache_if[i].req_data;
					// Trace: src/VX_cache_wrap.sv:86:5
					assign mem_bus_cache_if[i].req_ready = mem_bus_tmp_if[i].req_ready;
					// Trace: src/VX_cache_wrap.sv:87:5
					assign mem_bus_cache_if[i].rsp_valid = mem_bus_tmp_if[i].rsp_valid;
					// Trace: src/VX_cache_wrap.sv:88:5
					assign mem_bus_cache_if[i].rsp_data = mem_bus_tmp_if[i].rsp_data;
					// Trace: src/VX_cache_wrap.sv:89:5
					assign mem_bus_tmp_if[i].rsp_ready = mem_bus_cache_if[i].rsp_ready;
				end
			end
			// Trace: src/VX_cache_wrap.sv:92:5
			genvar _gv_i_169;
			for (_gv_i_169 = 0; _gv_i_169 < MEM_PORTS; _gv_i_169 = _gv_i_169 + 1) begin : g_mem_bus_if
				localparam i = _gv_i_169;
				if (WRITE_ENABLE) begin : g_we
					// Trace: src/VX_cache_wrap.sv:94:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
					// Trace: src/VX_cache_wrap.sv:95:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
					// Trace: src/VX_cache_wrap.sv:96:5
					assign mem_bus_tmp_if[i].req_ready = Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_ready;
					// Trace: src/VX_cache_wrap.sv:97:5
					assign mem_bus_tmp_if[i].rsp_valid = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
					// Trace: src/VX_cache_wrap.sv:98:5
					assign mem_bus_tmp_if[i].rsp_data = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
					// Trace: src/VX_cache_wrap.sv:99:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
				end
				else begin : g_ro
					// Trace: src/VX_cache_wrap.sv:101:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
					// Trace: src/VX_cache_wrap.sv:102:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[612] = 0;
					// Trace: src/VX_cache_wrap.sv:103:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[611-:26] = mem_bus_tmp_if[i].req_data[538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))-:((602 + (_param_4FE36_TAG_WIDTH + 2)) >= (579 + (_param_4FE36_TAG_WIDTH + 0)) ? ((538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))) - (512 + (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0))))) + 1 : ((512 + (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0)))) - (538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)))) + 1)];
					// Trace: src/VX_cache_wrap.sv:104:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[585-:512] = 1'sb0;
					// Trace: src/VX_cache_wrap.sv:105:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[73-:64] = 1'sb1;
					// Trace: src/VX_cache_wrap.sv:106:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[9-:3] = mem_bus_tmp_if[i].req_data[_param_4FE36_TAG_WIDTH + 2-:((_param_4FE36_TAG_WIDTH + 2) >= (_param_4FE36_TAG_WIDTH + 0) ? ((_param_4FE36_TAG_WIDTH + 2) - (_param_4FE36_TAG_WIDTH + 0)) + 1 : ((_param_4FE36_TAG_WIDTH + 0) - (_param_4FE36_TAG_WIDTH + 2)) + 1)];
					// Trace: src/VX_cache_wrap.sv:107:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[6-:7] = mem_bus_tmp_if[i].req_data[_param_4FE36_TAG_WIDTH - 1-:_param_4FE36_TAG_WIDTH + 0];
					// Trace: src/VX_cache_wrap.sv:108:5
					assign mem_bus_tmp_if[i].req_ready = Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_ready;
					// Trace: src/VX_cache_wrap.sv:109:5
					assign mem_bus_tmp_if[i].rsp_valid = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
					// Trace: src/VX_cache_wrap.sv:110:5
					assign mem_bus_tmp_if[i].rsp_data[_param_4FE36_TAG_WIDTH + 511-:((_param_4FE36_TAG_WIDTH + 511) >= (_param_4FE36_TAG_WIDTH + 0) ? ((_param_4FE36_TAG_WIDTH + 511) - (_param_4FE36_TAG_WIDTH + 0)) + 1 : ((_param_4FE36_TAG_WIDTH + 0) - (_param_4FE36_TAG_WIDTH + 511)) + 1)] = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_data[518-:512];
					// Trace: src/VX_cache_wrap.sv:111:5
					assign mem_bus_tmp_if[i].rsp_data[_param_4FE36_TAG_WIDTH - 1-:_param_4FE36_TAG_WIDTH + 0] = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_data[6-:7];
					// Trace: src/VX_cache_wrap.sv:112:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
				end
			end
			// Trace: src/VX_cache_wrap.sv:115:5
			if (1) begin : g_passthru
				genvar _gv_i_170;
				for (_gv_i_170 = 0; _gv_i_170 < NUM_REQS; _gv_i_170 = _gv_i_170 + 1) begin : g_core_bus_cache_if
					localparam i = _gv_i_170;
					// Trace: src/VX_cache_wrap.sv:146:5
					assign core_bus_cache_if[i].req_ready = 0;
					// Trace: src/VX_cache_wrap.sv:147:5
					assign core_bus_cache_if[i].rsp_valid = 0;
					// Trace: src/VX_cache_wrap.sv:148:5
					assign core_bus_cache_if[i].rsp_data = 1'sb0;
				end
				genvar _gv_i_171;
				for (_gv_i_171 = 0; _gv_i_171 < MEM_PORTS; _gv_i_171 = _gv_i_171 + 1) begin : g_mem_bus_cache_if
					localparam i = _gv_i_171;
					// Trace: src/VX_cache_wrap.sv:151:5
					assign mem_bus_cache_if[i].req_valid = 0;
					// Trace: src/VX_cache_wrap.sv:152:5
					assign mem_bus_cache_if[i].req_data = 1'sb0;
					// Trace: src/VX_cache_wrap.sv:153:5
					assign mem_bus_cache_if[i].rsp_ready = 0;
				end
			end
		end
	endgenerate
	assign l3cache.clk = clk;
	assign l3cache.reset = l3_reset;
	// Trace: src/Vortex.sv:64:5
	genvar _gv_i_123;
	generate
		for (_gv_i_123 = 0; _gv_i_123 < VX_gpu_pkg_L3_NUM_REQS; _gv_i_123 = _gv_i_123 + 1) begin : g_mem_bus_if
			localparam i = _gv_i_123;
			// Trace: src/Vortex.sv:65:9
			assign mem_req_valid[i] = mem_bus_if[i].req_valid;
			// Trace: src/Vortex.sv:66:9
			assign mem_req_rw[i] = mem_bus_if[i].req_data[612];
			// Trace: src/Vortex.sv:67:9
			assign mem_req_byteen[i * 64+:64] = mem_bus_if[i].req_data[73-:64];
			// Trace: src/Vortex.sv:68:9
			assign mem_req_addr[i * 26+:26] = mem_bus_if[i].req_data[611-:26];
			// Trace: src/Vortex.sv:69:9
			assign mem_req_data[i * 512+:512] = mem_bus_if[i].req_data[585-:512];
			// Trace: src/Vortex.sv:70:9
			assign mem_req_tag[i * 7+:7] = mem_bus_if[i].req_data[6-:7];
			// Trace: src/Vortex.sv:71:9
			assign mem_bus_if[i].req_ready = mem_req_ready[i];
			// Trace: src/Vortex.sv:72:9
			assign mem_bus_if[i].rsp_valid = mem_rsp_valid[i];
			// Trace: src/Vortex.sv:73:9
			assign mem_bus_if[i].rsp_data[518-:512] = mem_rsp_data[i * 512+:512];
			// Trace: src/Vortex.sv:74:9
			assign mem_bus_if[i].rsp_data[6-:7] = mem_rsp_tag[i * 7+:7];
			// Trace: src/Vortex.sv:75:9
			assign mem_rsp_ready[i] = mem_bus_if[i].rsp_ready;
		end
	endgenerate
	// Trace: src/Vortex.sv:77:5
	// expanded interface instance: dcr_bus_if
	generate
		if (1) begin : dcr_bus_if
			// Trace: src/VX_dcr_bus_if.sv:2:5
			wire write_valid;
			// Trace: src/VX_dcr_bus_if.sv:3:5
			wire [11:0] write_addr;
			// Trace: src/VX_dcr_bus_if.sv:4:5
			wire [31:0] write_data;
			// Trace: src/VX_dcr_bus_if.sv:5:5
			// Trace: src/VX_dcr_bus_if.sv:10:5
		end
	endgenerate
	// Trace: src/Vortex.sv:78:5
	assign dcr_bus_if.write_valid = dcr_wr_valid;
	// Trace: src/Vortex.sv:79:5
	assign dcr_bus_if.write_addr = dcr_wr_addr;
	// Trace: src/Vortex.sv:80:5
	assign dcr_bus_if.write_data = dcr_wr_data;
	// Trace: src/Vortex.sv:81:5
	wire [0:0] per_cluster_busy;
	// Trace: src/Vortex.sv:82:5
	genvar _gv_cluster_id_1;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	function automatic signed [2:0] sv2v_cast_22555_signed;
		input reg signed [2:0] inp;
		sv2v_cast_22555_signed = inp;
	endfunction
	function automatic signed [1:0] sv2v_cast_2_signed;
		input reg signed [1:0] inp;
		sv2v_cast_2_signed = inp;
	endfunction
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	function automatic signed [2:0] sv2v_cast_3_signed;
		input reg signed [2:0] inp;
		sv2v_cast_3_signed = inp;
	endfunction
	function automatic signed [0:0] sv2v_cast_1_signed;
		input reg signed [0:0] inp;
		sv2v_cast_1_signed = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [25:0] sv2v_cast_26;
		input reg [25:0] inp;
		sv2v_cast_26 = inp;
	endfunction
	function automatic signed [1:0] sv2v_cast_2C231_signed;
		input reg signed [1:0] inp;
		sv2v_cast_2C231_signed = inp;
	endfunction
	function automatic [43:0] sv2v_cast_44;
		input reg [43:0] inp;
		sv2v_cast_44 = inp;
	endfunction
	generate
		for (_gv_cluster_id_1 = 0; _gv_cluster_id_1 < 1; _gv_cluster_id_1 = _gv_cluster_id_1 + 1) begin : g_clusters
			localparam cluster_id = _gv_cluster_id_1;
			// Trace: src/Vortex.sv:83:5
			wire [0:0] cluster_reset;
			// Trace: src/Vortex.sv:84:5
			VX_reset_relay #(
				.N(1),
				.MAX_FANOUT(0)
			) __cluster_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(cluster_reset)
			);
			// Trace: src/Vortex.sv:89:9
			// expanded interface instance: cluster_dcr_bus_if
			if (1) begin : cluster_dcr_bus_if
				// Trace: src/VX_dcr_bus_if.sv:2:5
				wire write_valid;
				// Trace: src/VX_dcr_bus_if.sv:3:5
				wire [11:0] write_addr;
				// Trace: src/VX_dcr_bus_if.sv:4:5
				wire [31:0] write_data;
				// Trace: src/VX_dcr_bus_if.sv:5:5
				// Trace: src/VX_dcr_bus_if.sv:10:5
			end
			if (1) begin : genblk1
				// Trace: src/Vortex.sv:103:9
				assign {cluster_dcr_bus_if.write_valid, cluster_dcr_bus_if.write_addr, cluster_dcr_bus_if.write_data} = {dcr_bus_if.write_valid && 1'b1, dcr_bus_if.write_addr, dcr_bus_if.write_data};
			end
			// Trace: src/Vortex.sv:106:9
			// expanded module instance: cluster
			localparam _bbase_5867A_mem_bus_if = cluster_id * VX_gpu_pkg_L2_NUM_REQS;
			localparam _param_5867A_CLUSTER_ID = cluster_id;
			localparam _param_5867A_INSTANCE_ID = "";
			if (1) begin : cluster
				// removed import VX_gpu_pkg::*;
				// Trace: src/VX_cluster.sv:2:15
				localparam CLUSTER_ID = _param_5867A_CLUSTER_ID;
				// Trace: src/VX_cluster.sv:3:16
				localparam INSTANCE_ID = _param_5867A_INSTANCE_ID;
				// Trace: src/VX_cluster.sv:5:5
				wire clk;
				// Trace: src/VX_cluster.sv:6:5
				wire reset;
				// Trace: src/VX_cluster.sv:7:5
				// removed modport instance dcr_bus_if
				// Trace: src/VX_cluster.sv:8:5
				localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
				localparam VX_gpu_pkg_LSU_WORD_SIZE = 4;
				localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
				localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
				localparam VX_gpu_pkg_L2_NUM_REQS = 1;
				localparam _mbase_mem_bus_if = _bbase_5867A_mem_bus_if;
				// Trace: src/VX_cluster.sv:9:5
				wire busy;
				// Trace: src/VX_cluster.sv:11:5
				localparam VX_gpu_pkg_DCACHE_LINE_SIZE = 64;
				localparam VX_gpu_pkg_DCACHE_MERGED_REQS = 1;
				localparam VX_gpu_pkg_DCACHE_MEM_BATCHES = 1;
				localparam VX_gpu_pkg_DCACHE_TAG_ID_BITS = 2;
				localparam VX_gpu_pkg_DCACHE_TAG_WIDTH = 3;
				localparam VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH = 6;
				localparam VX_gpu_pkg_ICACHE_MEM_TAG_WIDTH = 5;
				localparam VX_gpu_pkg_L1_MEM_TAG_WIDTH = VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH;
				localparam VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH = 7;
				// expanded interface instance: per_socket_mem_bus_if
				localparam _param_1BD2B_DATA_SIZE = 64;
				localparam _param_1BD2B_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
				genvar _arr_1BD2B;
				for (_arr_1BD2B = 0; _arr_1BD2B <= 0; _arr_1BD2B = _arr_1BD2B + 1) begin : per_socket_mem_bus_if
					// Trace: src/VX_mem_bus_if.sv:2:15
					localparam DATA_SIZE = _param_1BD2B_DATA_SIZE;
					// Trace: src/VX_mem_bus_if.sv:3:15
					localparam FLAGS_WIDTH = 3;
					// Trace: src/VX_mem_bus_if.sv:4:15
					localparam TAG_WIDTH = _param_1BD2B_TAG_WIDTH;
					// Trace: src/VX_mem_bus_if.sv:5:15
					localparam MEM_ADDR_WIDTH = 32;
					// Trace: src/VX_mem_bus_if.sv:6:15
					localparam ADDR_WIDTH = 26;
					// Trace: src/VX_mem_bus_if.sv:7:15
					localparam UUID_WIDTH = 1;
					// Trace: src/VX_mem_bus_if.sv:9:5
					// removed localparam type tag_t
					// Trace: src/VX_mem_bus_if.sv:13:5
					// removed localparam type req_data_t
					// Trace: src/VX_mem_bus_if.sv:21:5
					// removed localparam type rsp_data_t
					// Trace: src/VX_mem_bus_if.sv:25:5
					wire req_valid;
					// Trace: src/VX_mem_bus_if.sv:26:5
					wire [612:0] req_data;
					// Trace: src/VX_mem_bus_if.sv:27:5
					wire req_ready;
					// Trace: src/VX_mem_bus_if.sv:28:5
					wire rsp_valid;
					// Trace: src/VX_mem_bus_if.sv:29:5
					wire [518:0] rsp_data;
					// Trace: src/VX_mem_bus_if.sv:30:5
					wire rsp_ready;
					// Trace: src/VX_mem_bus_if.sv:31:5
					// Trace: src/VX_mem_bus_if.sv:39:5
				end
				// Trace: src/VX_cluster.sv:15:5
				wire [0:0] l2_reset;
				// Trace: src/VX_cluster.sv:16:5
				VX_reset_relay #(
					.N(1),
					.MAX_FANOUT(0)
				) __l2_reset(
					.clk(clk),
					.reset(reset),
					.reset_o(l2_reset)
				);
				// Trace: src/VX_cluster.sv:21:5
				localparam VX_gpu_pkg_L2_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
				localparam VX_gpu_pkg_L2_WORD_SIZE = 64;
				// expanded module instance: l2cache
				localparam _bbase_56EB4_core_bus_if = 0;
				localparam _bbase_56EB4_mem_bus_if = cluster_id * VX_gpu_pkg_L2_NUM_REQS;
				localparam _param_56EB4_INSTANCE_ID = "";
				localparam _param_56EB4_CACHE_SIZE = 1048576;
				localparam _param_56EB4_LINE_SIZE = 64;
				localparam _param_56EB4_NUM_BANKS = VX_gpu_pkg_L2_NUM_REQS;
				localparam _param_56EB4_NUM_WAYS = 8;
				localparam _param_56EB4_WORD_SIZE = VX_gpu_pkg_L2_WORD_SIZE;
				localparam _param_56EB4_NUM_REQS = VX_gpu_pkg_L2_NUM_REQS;
				localparam _param_56EB4_MEM_PORTS = VX_gpu_pkg_L2_NUM_REQS;
				localparam _param_56EB4_CRSQ_SIZE = 2;
				localparam _param_56EB4_MSHR_SIZE = 16;
				localparam _param_56EB4_MRSQ_SIZE = 4;
				localparam _param_56EB4_MREQ_SIZE = 4;
				localparam _param_56EB4_TAG_WIDTH = VX_gpu_pkg_L2_TAG_WIDTH;
				localparam _param_56EB4_WRITE_ENABLE = 1;
				localparam _param_56EB4_WRITEBACK = 0;
				localparam _param_56EB4_DIRTY_BYTES = 0;
				localparam _param_56EB4_REPL_POLICY = 1;
				localparam _param_56EB4_UUID_WIDTH = 1;
				localparam _param_56EB4_FLAGS_WIDTH = 3;
				localparam _param_56EB4_CORE_OUT_BUF = 3;
				localparam _param_56EB4_MEM_OUT_BUF = 3;
				localparam _param_56EB4_NC_ENABLE = 1;
				localparam _param_56EB4_PASSTHRU = 1'd1;
				if (1) begin : l2cache
					// removed import VX_gpu_pkg::*;
					// Trace: src/VX_cache_wrap.sv:2:16
					localparam INSTANCE_ID = _param_56EB4_INSTANCE_ID;
					// Trace: src/VX_cache_wrap.sv:3:15
					localparam TAG_SEL_IDX = 0;
					// Trace: src/VX_cache_wrap.sv:4:15
					localparam NUM_REQS = _param_56EB4_NUM_REQS;
					// Trace: src/VX_cache_wrap.sv:5:15
					localparam MEM_PORTS = _param_56EB4_MEM_PORTS;
					// Trace: src/VX_cache_wrap.sv:6:15
					localparam CACHE_SIZE = _param_56EB4_CACHE_SIZE;
					// Trace: src/VX_cache_wrap.sv:7:15
					localparam LINE_SIZE = _param_56EB4_LINE_SIZE;
					// Trace: src/VX_cache_wrap.sv:8:15
					localparam NUM_BANKS = _param_56EB4_NUM_BANKS;
					// Trace: src/VX_cache_wrap.sv:9:15
					localparam NUM_WAYS = _param_56EB4_NUM_WAYS;
					// Trace: src/VX_cache_wrap.sv:10:15
					localparam WORD_SIZE = _param_56EB4_WORD_SIZE;
					// Trace: src/VX_cache_wrap.sv:11:15
					localparam CRSQ_SIZE = _param_56EB4_CRSQ_SIZE;
					// Trace: src/VX_cache_wrap.sv:12:15
					localparam MSHR_SIZE = _param_56EB4_MSHR_SIZE;
					// Trace: src/VX_cache_wrap.sv:13:15
					localparam MRSQ_SIZE = _param_56EB4_MRSQ_SIZE;
					// Trace: src/VX_cache_wrap.sv:14:15
					localparam MREQ_SIZE = _param_56EB4_MREQ_SIZE;
					// Trace: src/VX_cache_wrap.sv:15:15
					localparam WRITE_ENABLE = _param_56EB4_WRITE_ENABLE;
					// Trace: src/VX_cache_wrap.sv:16:15
					localparam WRITEBACK = _param_56EB4_WRITEBACK;
					// Trace: src/VX_cache_wrap.sv:17:15
					localparam DIRTY_BYTES = _param_56EB4_DIRTY_BYTES;
					// Trace: src/VX_cache_wrap.sv:18:15
					localparam REPL_POLICY = _param_56EB4_REPL_POLICY;
					// Trace: src/VX_cache_wrap.sv:19:15
					localparam UUID_WIDTH = _param_56EB4_UUID_WIDTH;
					// Trace: src/VX_cache_wrap.sv:20:15
					localparam TAG_WIDTH = _param_56EB4_TAG_WIDTH;
					// Trace: src/VX_cache_wrap.sv:21:15
					localparam FLAGS_WIDTH = _param_56EB4_FLAGS_WIDTH;
					// Trace: src/VX_cache_wrap.sv:22:15
					localparam NC_ENABLE = _param_56EB4_NC_ENABLE;
					// Trace: src/VX_cache_wrap.sv:23:15
					localparam PASSTHRU = _param_56EB4_PASSTHRU;
					// Trace: src/VX_cache_wrap.sv:24:15
					localparam CORE_OUT_BUF = _param_56EB4_CORE_OUT_BUF;
					// Trace: src/VX_cache_wrap.sv:25:15
					localparam MEM_OUT_BUF = _param_56EB4_MEM_OUT_BUF;
					// Trace: src/VX_cache_wrap.sv:27:5
					wire clk;
					// Trace: src/VX_cache_wrap.sv:28:5
					wire reset;
					// Trace: src/VX_cache_wrap.sv:29:5
					localparam _mbase_core_bus_if = 0;
					// Trace: src/VX_cache_wrap.sv:30:5
					localparam _mbase_mem_bus_if = _bbase_56EB4_mem_bus_if;
					// Trace: src/VX_cache_wrap.sv:32:5
					localparam CACHE_MEM_TAG_WIDTH = 5;
					// Trace: src/VX_cache_wrap.sv:34:5
					localparam BYPASS_TAG_WIDTH = 7;
					// Trace: src/VX_cache_wrap.sv:36:5
					localparam NC_TAG_WIDTH = 8;
					// Trace: src/VX_cache_wrap.sv:37:5
					localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
					// Trace: src/VX_cache_wrap.sv:38:5
					localparam BYPASS_ENABLE = 1'd1;
					// Trace: src/VX_cache_wrap.sv:39:5
					// expanded interface instance: core_bus_cache_if
					localparam _param_24C1C_DATA_SIZE = WORD_SIZE;
					localparam _param_24C1C_TAG_WIDTH = TAG_WIDTH;
					genvar _arr_24C1C;
					for (_arr_24C1C = 0; _arr_24C1C <= 0; _arr_24C1C = _arr_24C1C + 1) begin : core_bus_cache_if
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_24C1C_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_24C1C_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:7:15
						localparam UUID_WIDTH = 1;
						// Trace: src/VX_mem_bus_if.sv:9:5
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:13:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:21:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:30:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:31:5
						// Trace: src/VX_mem_bus_if.sv:39:5
					end
					// Trace: src/VX_cache_wrap.sv:43:5
					// expanded interface instance: mem_bus_cache_if
					localparam _param_D895D_DATA_SIZE = LINE_SIZE;
					localparam _param_D895D_TAG_WIDTH = CACHE_MEM_TAG_WIDTH;
					genvar _arr_D895D;
					for (_arr_D895D = 0; _arr_D895D <= 0; _arr_D895D = _arr_D895D + 1) begin : mem_bus_cache_if
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_D895D_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_D895D_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:7:15
						localparam UUID_WIDTH = 1;
						// Trace: src/VX_mem_bus_if.sv:9:5
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:13:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:21:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire [610:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire [516:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:30:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:31:5
						// Trace: src/VX_mem_bus_if.sv:39:5
					end
					// Trace: src/VX_cache_wrap.sv:47:5
					// expanded interface instance: mem_bus_tmp_if
					localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
					localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
					genvar _arr_4FE36;
					for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam FLAGS_WIDTH = 3;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:7:15
						localparam UUID_WIDTH = 1;
						// Trace: src/VX_mem_bus_if.sv:9:5
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:13:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:21:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:30:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:31:5
						// Trace: src/VX_mem_bus_if.sv:39:5
					end
					// Trace: src/VX_cache_wrap.sv:51:5
					if (BYPASS_ENABLE) begin : g_bypass
						// Trace: src/VX_cache_wrap.sv:52:9
						// expanded module instance: cache_bypass
						localparam _bbase_714AA_core_bus_in_if = 0;
						localparam _bbase_714AA_core_bus_out_if = 0;
						localparam _bbase_714AA_mem_bus_in_if = 0;
						localparam _bbase_714AA_mem_bus_out_if = 0;
						localparam _param_714AA_NUM_REQS = NUM_REQS;
						localparam _param_714AA_MEM_PORTS = MEM_PORTS;
						localparam _param_714AA_TAG_SEL_IDX = TAG_SEL_IDX;
						localparam _param_714AA_CACHE_ENABLE = !PASSTHRU;
						localparam _param_714AA_WORD_SIZE = WORD_SIZE;
						localparam _param_714AA_LINE_SIZE = LINE_SIZE;
						localparam _param_714AA_CORE_ADDR_WIDTH = 26;
						localparam _param_714AA_CORE_TAG_WIDTH = TAG_WIDTH;
						localparam _param_714AA_MEM_ADDR_WIDTH = 26;
						localparam _param_714AA_MEM_TAG_IN_WIDTH = CACHE_MEM_TAG_WIDTH;
						localparam _param_714AA_UUID_WIDTH = UUID_WIDTH;
						localparam _param_714AA_CORE_OUT_BUF = CORE_OUT_BUF;
						localparam _param_714AA_MEM_OUT_BUF = MEM_OUT_BUF;
						if (1) begin : cache_bypass
							// Trace: src/VX_cache_bypass.sv:2:15
							localparam NUM_REQS = _param_714AA_NUM_REQS;
							// Trace: src/VX_cache_bypass.sv:3:15
							localparam MEM_PORTS = _param_714AA_MEM_PORTS;
							// Trace: src/VX_cache_bypass.sv:4:15
							localparam TAG_SEL_IDX = _param_714AA_TAG_SEL_IDX;
							// Trace: src/VX_cache_bypass.sv:5:15
							localparam CACHE_ENABLE = _param_714AA_CACHE_ENABLE;
							// Trace: src/VX_cache_bypass.sv:6:15
							localparam WORD_SIZE = _param_714AA_WORD_SIZE;
							// Trace: src/VX_cache_bypass.sv:7:15
							localparam LINE_SIZE = _param_714AA_LINE_SIZE;
							// Trace: src/VX_cache_bypass.sv:8:15
							localparam CORE_ADDR_WIDTH = _param_714AA_CORE_ADDR_WIDTH;
							// Trace: src/VX_cache_bypass.sv:9:15
							localparam CORE_TAG_WIDTH = _param_714AA_CORE_TAG_WIDTH;
							// Trace: src/VX_cache_bypass.sv:10:15
							localparam MEM_ADDR_WIDTH = _param_714AA_MEM_ADDR_WIDTH;
							// Trace: src/VX_cache_bypass.sv:11:15
							localparam MEM_TAG_IN_WIDTH = _param_714AA_MEM_TAG_IN_WIDTH;
							// Trace: src/VX_cache_bypass.sv:12:15
							localparam UUID_WIDTH = _param_714AA_UUID_WIDTH;
							// Trace: src/VX_cache_bypass.sv:13:15
							localparam CORE_OUT_BUF = _param_714AA_CORE_OUT_BUF;
							// Trace: src/VX_cache_bypass.sv:14:15
							localparam MEM_OUT_BUF = _param_714AA_MEM_OUT_BUF;
							// Trace: src/VX_cache_bypass.sv:16:5
							wire clk;
							// Trace: src/VX_cache_bypass.sv:17:5
							wire reset;
							// Trace: src/VX_cache_bypass.sv:18:5
							localparam _mbase_core_bus_in_if = 0;
							// Trace: src/VX_cache_bypass.sv:19:5
							localparam _mbase_core_bus_out_if = 0;
							// Trace: src/VX_cache_bypass.sv:20:5
							localparam _mbase_mem_bus_in_if = 0;
							// Trace: src/VX_cache_bypass.sv:21:5
							localparam _mbase_mem_bus_out_if = 0;
							// Trace: src/VX_cache_bypass.sv:23:5
							localparam DIRECT_PASSTHRU = (!CACHE_ENABLE && 1'd1) && 1'd1;
							// Trace: src/VX_cache_bypass.sv:24:5
							localparam CORE_DATA_WIDTH = 512;
							// Trace: src/VX_cache_bypass.sv:25:5
							localparam WORDS_PER_LINE = 1;
							// Trace: src/VX_cache_bypass.sv:26:5
							localparam WSEL_BITS = 0;
							// Trace: src/VX_cache_bypass.sv:27:5
							localparam CORE_TAG_ID_WIDTH = 6;
							// Trace: src/VX_cache_bypass.sv:28:5
							localparam MEM_TAG_ID_WIDTH = 6;
							// Trace: src/VX_cache_bypass.sv:29:5
							localparam MEM_TAG_NC1_WIDTH = 7;
							// Trace: src/VX_cache_bypass.sv:30:5
							localparam MEM_TAG_NC2_WIDTH = 7;
							// Trace: src/VX_cache_bypass.sv:31:5
							localparam MEM_TAG_OUT_WIDTH = (CACHE_ENABLE ? MEM_TAG_NC2_WIDTH : MEM_TAG_NC2_WIDTH);
							// Trace: src/VX_cache_bypass.sv:32:5
							// expanded interface instance: core_bus_nc_switch_if
							localparam _param_95306_DATA_SIZE = WORD_SIZE;
							localparam _param_95306_TAG_WIDTH = CORE_TAG_WIDTH;
							genvar _arr_95306;
							for (_arr_95306 = 0; _arr_95306 <= (((CACHE_ENABLE ? 2 : 1) * NUM_REQS) - 1); _arr_95306 = _arr_95306 + 1) begin : core_bus_nc_switch_if
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_95306_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_95306_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:7:15
								localparam UUID_WIDTH = 1;
								// Trace: src/VX_mem_bus_if.sv:9:5
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:13:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:21:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:30:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:31:5
								// Trace: src/VX_mem_bus_if.sv:39:5
							end
							// Trace: src/VX_cache_bypass.sv:36:5
							wire [0:0] core_req_nc_sel;
							// Trace: src/VX_cache_bypass.sv:37:5
							genvar _gv_i_179;
							for (_gv_i_179 = 0; _gv_i_179 < NUM_REQS; _gv_i_179 = _gv_i_179 + 1) begin : g_core_req_is_nc
								localparam i = _gv_i_179;
								if (CACHE_ENABLE) begin : g_cache
									// Trace: src/VX_cache_bypass.sv:39:13
									assign core_req_nc_sel[i] = ~Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_in_if].req_data[8];
								end
								else begin : g_no_cache
									// Trace: src/VX_cache_bypass.sv:41:13
									assign core_req_nc_sel[i] = 1'b0;
								end
							end
							// Trace: src/VX_cache_bypass.sv:44:5
							// expanded module instance: core_bus_nc_switch
							localparam _bbase_69FDB_bus_in_if = 0;
							localparam _bbase_69FDB_bus_out_if = 0;
							localparam _param_69FDB_NUM_INPUTS = NUM_REQS;
							localparam _param_69FDB_NUM_OUTPUTS = (CACHE_ENABLE ? 2 : 1) * NUM_REQS;
							localparam _param_69FDB_DATA_SIZE = WORD_SIZE;
							localparam _param_69FDB_TAG_WIDTH = CORE_TAG_WIDTH;
							localparam _param_69FDB_ARBITER = "R";
							localparam _param_69FDB_REQ_OUT_BUF = 0;
							localparam _param_69FDB_RSP_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
							if (1) begin : core_bus_nc_switch
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_switch.sv:2:15
								localparam NUM_INPUTS = _param_69FDB_NUM_INPUTS;
								// Trace: src/VX_mem_switch.sv:3:15
								localparam NUM_OUTPUTS = _param_69FDB_NUM_OUTPUTS;
								// Trace: src/VX_mem_switch.sv:4:15
								localparam DATA_SIZE = _param_69FDB_DATA_SIZE;
								// Trace: src/VX_mem_switch.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_switch.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_switch.sv:7:15
								localparam TAG_WIDTH = _param_69FDB_TAG_WIDTH;
								// Trace: src/VX_mem_switch.sv:8:15
								localparam REQ_OUT_BUF = _param_69FDB_REQ_OUT_BUF;
								// Trace: src/VX_mem_switch.sv:9:15
								localparam RSP_OUT_BUF = _param_69FDB_RSP_OUT_BUF;
								// Trace: src/VX_mem_switch.sv:10:16
								localparam ARBITER = _param_69FDB_ARBITER;
								// Trace: src/VX_mem_switch.sv:11:15
								localparam NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
								// Trace: src/VX_mem_switch.sv:12:15
								localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
								// Trace: src/VX_mem_switch.sv:13:15
								localparam LOG_NUM_REQS = $clog2(NUM_REQS);
								// Trace: src/VX_mem_switch.sv:15:5
								wire clk;
								// Trace: src/VX_mem_switch.sv:16:5
								wire reset;
								// Trace: src/VX_mem_switch.sv:17:5
								wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] bus_sel;
								// Trace: src/VX_mem_switch.sv:18:5
								localparam _mbase_bus_in_if = 0;
								// Trace: src/VX_mem_switch.sv:19:5
								localparam _mbase_bus_out_if = 0;
								// Trace: src/VX_mem_switch.sv:21:5
								localparam DATA_WIDTH = 512;
								// Trace: src/VX_mem_switch.sv:22:5
								localparam REQ_DATAW = 613;
								// Trace: src/VX_mem_switch.sv:23:5
								localparam RSP_DATAW = 519;
								// Trace: src/VX_mem_switch.sv:24:5
								wire [0:0] req_valid_in;
								// Trace: src/VX_mem_switch.sv:25:5
								wire [612:0] req_data_in;
								// Trace: src/VX_mem_switch.sv:26:5
								wire [0:0] req_ready_in;
								// Trace: src/VX_mem_switch.sv:27:5
								wire [NUM_OUTPUTS - 1:0] req_valid_out;
								// Trace: src/VX_mem_switch.sv:28:5
								wire [(NUM_OUTPUTS * 613) - 1:0] req_data_out;
								// Trace: src/VX_mem_switch.sv:29:5
								wire [NUM_OUTPUTS - 1:0] req_ready_out;
								// Trace: src/VX_mem_switch.sv:30:5
								genvar _gv_i_154;
								for (_gv_i_154 = 0; _gv_i_154 < NUM_INPUTS; _gv_i_154 = _gv_i_154 + 1) begin : g_req_data_in
									localparam i = _gv_i_154;
									// Trace: src/VX_mem_switch.sv:31:9
									assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].req_valid;
									// Trace: src/VX_mem_switch.sv:32:9
									assign req_data_in[i * 613+:613] = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].req_data;
									// Trace: src/VX_mem_switch.sv:33:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
								end
								// Trace: src/VX_mem_switch.sv:35:5
								VX_stream_switch #(
									.NUM_INPUTS(NUM_INPUTS),
									.NUM_OUTPUTS(NUM_OUTPUTS),
									.DATAW(REQ_DATAW),
									.OUT_BUF(REQ_OUT_BUF)
								) req_switch(
									.clk(clk),
									.reset(reset),
									.sel_in(bus_sel),
									.valid_in(req_valid_in),
									.data_in(req_data_in),
									.ready_in(req_ready_in),
									.valid_out(req_valid_out),
									.data_out(req_data_out),
									.ready_out(req_ready_out)
								);
								// Trace: src/VX_mem_switch.sv:51:5
								genvar _gv_i_155;
								for (_gv_i_155 = 0; _gv_i_155 < NUM_OUTPUTS; _gv_i_155 = _gv_i_155 + 1) begin : g_req_data_out
									localparam i = _gv_i_155;
									// Trace: src/VX_mem_switch.sv:52:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
									// Trace: src/VX_mem_switch.sv:53:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_data = req_data_out[i * 613+:613];
									// Trace: src/VX_mem_switch.sv:54:9
									assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_ready;
								end
								// Trace: src/VX_mem_switch.sv:56:5
								wire [NUM_OUTPUTS - 1:0] rsp_valid_in;
								// Trace: src/VX_mem_switch.sv:57:5
								wire [(NUM_OUTPUTS * 519) - 1:0] rsp_data_in;
								// Trace: src/VX_mem_switch.sv:58:5
								wire [NUM_OUTPUTS - 1:0] rsp_ready_in;
								// Trace: src/VX_mem_switch.sv:59:5
								wire [0:0] rsp_valid_out;
								// Trace: src/VX_mem_switch.sv:60:5
								wire [518:0] rsp_data_out;
								// Trace: src/VX_mem_switch.sv:61:5
								wire [0:0] rsp_ready_out;
								// Trace: src/VX_mem_switch.sv:62:5
								genvar _gv_i_156;
								for (_gv_i_156 = 0; _gv_i_156 < NUM_OUTPUTS; _gv_i_156 = _gv_i_156 + 1) begin : g_rsp_data_in
									localparam i = _gv_i_156;
									// Trace: src/VX_mem_switch.sv:63:9
									assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_valid;
									// Trace: src/VX_mem_switch.sv:64:9
									assign rsp_data_in[i * 519+:519] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_data;
									// Trace: src/VX_mem_switch.sv:65:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
								end
								// Trace: src/VX_mem_switch.sv:67:5
								VX_stream_arb #(
									.NUM_INPUTS(NUM_OUTPUTS),
									.NUM_OUTPUTS(NUM_INPUTS),
									.DATAW(RSP_DATAW),
									.ARBITER(ARBITER),
									.OUT_BUF(RSP_OUT_BUF)
								) rsp_arb(
									.clk(clk),
									.reset(reset),
									.valid_in(rsp_valid_in),
									.data_in(rsp_data_in),
									.ready_in(rsp_ready_in),
									.valid_out(rsp_valid_out),
									.data_out(rsp_data_out),
									.ready_out(rsp_ready_out),
									.sel_out()
								);
								// Trace: src/VX_mem_switch.sv:84:5
								genvar _gv_i_157;
								for (_gv_i_157 = 0; _gv_i_157 < NUM_INPUTS; _gv_i_157 = _gv_i_157 + 1) begin : g_rsp_data_out
									localparam i = _gv_i_157;
									// Trace: src/VX_mem_switch.sv:85:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
									// Trace: src/VX_mem_switch.sv:86:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
									// Trace: src/VX_mem_switch.sv:87:9
									assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].rsp_ready;
								end
							end
							assign core_bus_nc_switch.clk = clk;
							assign core_bus_nc_switch.reset = reset;
							assign core_bus_nc_switch.bus_sel = core_req_nc_sel;
							// Trace: src/VX_cache_bypass.sv:59:5
							// expanded interface instance: core_bus_in_nc_if
							localparam _param_C0263_DATA_SIZE = WORD_SIZE;
							localparam _param_C0263_TAG_WIDTH = CORE_TAG_WIDTH;
							genvar _arr_C0263;
							for (_arr_C0263 = 0; _arr_C0263 <= 0; _arr_C0263 = _arr_C0263 + 1) begin : core_bus_in_nc_if
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_C0263_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_C0263_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:7:15
								localparam UUID_WIDTH = 1;
								// Trace: src/VX_mem_bus_if.sv:9:5
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:13:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:21:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:30:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:31:5
								// Trace: src/VX_mem_bus_if.sv:39:5
							end
							// Trace: src/VX_cache_bypass.sv:63:5
							genvar _gv_i_180;
							for (_gv_i_180 = 0; _gv_i_180 < NUM_REQS; _gv_i_180 = _gv_i_180 + 1) begin : g_core_bus_nc_switch_if
								localparam i = _gv_i_180;
								// Trace: src/VX_cache_bypass.sv:64:9
								assign core_bus_in_nc_if[i].req_valid = core_bus_nc_switch_if[0 + i].req_valid;
								// Trace: src/VX_cache_bypass.sv:65:9
								assign core_bus_in_nc_if[i].req_data = core_bus_nc_switch_if[0 + i].req_data;
								// Trace: src/VX_cache_bypass.sv:66:9
								assign core_bus_nc_switch_if[0 + i].req_ready = core_bus_in_nc_if[i].req_ready;
								// Trace: src/VX_cache_bypass.sv:67:9
								assign core_bus_nc_switch_if[0 + i].rsp_valid = core_bus_in_nc_if[i].rsp_valid;
								// Trace: src/VX_cache_bypass.sv:68:9
								assign core_bus_nc_switch_if[0 + i].rsp_data = core_bus_in_nc_if[i].rsp_data;
								// Trace: src/VX_cache_bypass.sv:69:9
								assign core_bus_in_nc_if[i].rsp_ready = core_bus_nc_switch_if[0 + i].rsp_ready;
								if (CACHE_ENABLE) begin : g_cache
									// Trace: src/VX_cache_bypass.sv:71:13
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = core_bus_nc_switch_if[1 + i].req_valid;
									// Trace: src/VX_cache_bypass.sv:72:13
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = core_bus_nc_switch_if[1 + i].req_data;
									// Trace: src/VX_cache_bypass.sv:73:13
									assign core_bus_nc_switch_if[1 + i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_ready;
									// Trace: src/VX_cache_bypass.sv:74:13
									assign core_bus_nc_switch_if[1 + i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_valid;
									// Trace: src/VX_cache_bypass.sv:75:13
									assign core_bus_nc_switch_if[1 + i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_data;
									// Trace: src/VX_cache_bypass.sv:76:13
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = core_bus_nc_switch_if[1 + i].rsp_ready;
								end
								else begin : g_no_cache
									// Trace: src/VX_cache_bypass.sv:78:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = 0;
									// Trace: src/VX_cache_bypass.sv:79:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = 1'sb0;
									// Trace: src/VX_cache_bypass.sv:80:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = 0;
								end
							end
							// Trace: src/VX_cache_bypass.sv:83:5
							// expanded interface instance: core_bus_nc_arb_if
							localparam _param_D50AC_DATA_SIZE = WORD_SIZE;
							localparam _param_D50AC_TAG_WIDTH = MEM_TAG_NC1_WIDTH;
							genvar _arr_D50AC;
							for (_arr_D50AC = 0; _arr_D50AC <= 0; _arr_D50AC = _arr_D50AC + 1) begin : core_bus_nc_arb_if
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_D50AC_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_D50AC_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:7:15
								localparam UUID_WIDTH = 1;
								// Trace: src/VX_mem_bus_if.sv:9:5
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:13:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:21:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:30:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:31:5
								// Trace: src/VX_mem_bus_if.sv:39:5
							end
							// Trace: src/VX_cache_bypass.sv:87:5
							// expanded module instance: core_bus_nc_arb
							localparam _bbase_1376F_bus_in_if = 0;
							localparam _bbase_1376F_bus_out_if = 0;
							localparam _param_1376F_NUM_INPUTS = NUM_REQS;
							localparam _param_1376F_NUM_OUTPUTS = MEM_PORTS;
							localparam _param_1376F_DATA_SIZE = WORD_SIZE;
							localparam _param_1376F_TAG_WIDTH = CORE_TAG_WIDTH;
							localparam _param_1376F_TAG_SEL_IDX = TAG_SEL_IDX;
							localparam _param_1376F_ARBITER = (CACHE_ENABLE ? "P" : "R");
							localparam _param_1376F_REQ_OUT_BUF = 0;
							localparam _param_1376F_RSP_OUT_BUF = 0;
							if (1) begin : core_bus_nc_arb
								// Trace: src/VX_mem_arb.sv:2:15
								localparam NUM_INPUTS = _param_1376F_NUM_INPUTS;
								// Trace: src/VX_mem_arb.sv:3:15
								localparam NUM_OUTPUTS = _param_1376F_NUM_OUTPUTS;
								// Trace: src/VX_mem_arb.sv:4:15
								localparam DATA_SIZE = _param_1376F_DATA_SIZE;
								// Trace: src/VX_mem_arb.sv:5:15
								localparam TAG_WIDTH = _param_1376F_TAG_WIDTH;
								// Trace: src/VX_mem_arb.sv:6:15
								localparam TAG_SEL_IDX = _param_1376F_TAG_SEL_IDX;
								// Trace: src/VX_mem_arb.sv:7:15
								localparam REQ_OUT_BUF = _param_1376F_REQ_OUT_BUF;
								// Trace: src/VX_mem_arb.sv:8:15
								localparam RSP_OUT_BUF = _param_1376F_RSP_OUT_BUF;
								// Trace: src/VX_mem_arb.sv:9:16
								localparam ARBITER = _param_1376F_ARBITER;
								// Trace: src/VX_mem_arb.sv:10:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_arb.sv:11:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_arb.sv:12:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_arb.sv:14:5
								wire clk;
								// Trace: src/VX_mem_arb.sv:15:5
								wire reset;
								// Trace: src/VX_mem_arb.sv:16:5
								localparam _mbase_bus_in_if = 0;
								// Trace: src/VX_mem_arb.sv:17:5
								localparam _mbase_bus_out_if = 0;
								// Trace: src/VX_mem_arb.sv:19:5
								localparam DATA_WIDTH = 512;
								// Trace: src/VX_mem_arb.sv:20:5
								localparam LOG_NUM_REQS = 0;
								// Trace: src/VX_mem_arb.sv:21:5
								localparam REQ_DATAW = 613;
								// Trace: src/VX_mem_arb.sv:22:5
								localparam RSP_DATAW = 519;
								// Trace: src/VX_mem_arb.sv:24:5
								wire [0:0] req_valid_in;
								// Trace: src/VX_mem_arb.sv:25:5
								wire [612:0] req_data_in;
								// Trace: src/VX_mem_arb.sv:26:5
								wire [0:0] req_ready_in;
								// Trace: src/VX_mem_arb.sv:27:5
								wire [0:0] req_valid_out;
								// Trace: src/VX_mem_arb.sv:28:5
								wire [612:0] req_data_out;
								// Trace: src/VX_mem_arb.sv:29:5
								wire [0:0] req_sel_out;
								// Trace: src/VX_mem_arb.sv:30:5
								wire [0:0] req_ready_out;
								// Trace: src/VX_mem_arb.sv:31:5
								genvar _gv_i_80;
								for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
									localparam i = _gv_i_80;
									// Trace: src/VX_mem_arb.sv:32:9
									assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_valid;
									// Trace: src/VX_mem_arb.sv:33:9
									assign req_data_in[i * 613+:613] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_data;
									// Trace: src/VX_mem_arb.sv:34:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
								end
								// Trace: src/VX_mem_arb.sv:36:5
								VX_stream_arb #(
									.NUM_INPUTS(NUM_INPUTS),
									.NUM_OUTPUTS(NUM_OUTPUTS),
									.DATAW(REQ_DATAW),
									.ARBITER(ARBITER),
									.OUT_BUF(REQ_OUT_BUF)
								) req_arb(
									.clk(clk),
									.reset(reset),
									.valid_in(req_valid_in),
									.ready_in(req_ready_in),
									.data_in(req_data_in),
									.data_out(req_data_out),
									.sel_out(req_sel_out),
									.valid_out(req_valid_out),
									.ready_out(req_ready_out)
								);
								// Trace: src/VX_mem_arb.sv:53:5
								genvar _gv_i_81;
								for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
									localparam i = _gv_i_81;
									// Trace: src/VX_mem_arb.sv:54:9
									wire [6:0] req_tag_out;
									// Trace: src/VX_mem_arb.sv:55:9
									VX_bits_insert #(
										.N(TAG_WIDTH),
										.S(LOG_NUM_REQS),
										.POS(TAG_SEL_IDX)
									) bits_insert(
										.data_in(req_tag_out),
										.ins_in(req_sel_out[i+:1]),
										.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[6-:7])
									);
									// Trace: src/VX_mem_arb.sv:64:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
									// Trace: src/VX_mem_arb.sv:65:9
									assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[612], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[611-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[585-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[73-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[9-:3], req_tag_out} = req_data_out[i * 613+:613];
									// Trace: src/VX_mem_arb.sv:73:9
									assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_ready;
								end
								// Trace: src/VX_mem_arb.sv:75:5
								wire [0:0] rsp_valid_out;
								// Trace: src/VX_mem_arb.sv:76:5
								wire [518:0] rsp_data_out;
								// Trace: src/VX_mem_arb.sv:77:5
								wire [0:0] rsp_ready_out;
								// Trace: src/VX_mem_arb.sv:78:5
								wire [0:0] rsp_valid_in;
								// Trace: src/VX_mem_arb.sv:79:5
								wire [518:0] rsp_data_in;
								// Trace: src/VX_mem_arb.sv:80:5
								wire [0:0] rsp_ready_in;
								// Trace: src/VX_mem_arb.sv:81:5
								if (1) begin : g_passthru
									genvar _gv_i_83;
									for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
										localparam i = _gv_i_83;
										// Trace: src/VX_mem_arb.sv:116:13
										assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_valid;
										// Trace: src/VX_mem_arb.sv:117:13
										assign rsp_data_in[i * 519+:519] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_data;
										// Trace: src/VX_mem_arb.sv:118:13
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:120:9
									VX_stream_arb #(
										.NUM_INPUTS(NUM_OUTPUTS),
										.NUM_OUTPUTS(NUM_INPUTS),
										.DATAW(RSP_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(RSP_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(rsp_valid_in),
										.ready_in(rsp_ready_in),
										.data_in(rsp_data_in),
										.data_out(rsp_data_out),
										.valid_out(rsp_valid_out),
										.ready_out(rsp_ready_out),
										.sel_out()
									);
								end
								// Trace: src/VX_mem_arb.sv:138:5
								genvar _gv_i_84;
								for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
									localparam i = _gv_i_84;
									// Trace: src/VX_mem_arb.sv:139:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
									// Trace: src/VX_mem_arb.sv:140:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
									// Trace: src/VX_mem_arb.sv:141:9
									assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_ready;
								end
							end
							assign core_bus_nc_arb.clk = clk;
							assign core_bus_nc_arb.reset = reset;
							// Trace: src/VX_cache_bypass.sv:102:5
							// expanded interface instance: mem_bus_out_nc_if
							localparam _param_0061C_DATA_SIZE = LINE_SIZE;
							localparam _param_0061C_TAG_WIDTH = MEM_TAG_NC2_WIDTH;
							genvar _arr_0061C;
							for (_arr_0061C = 0; _arr_0061C <= 0; _arr_0061C = _arr_0061C + 1) begin : mem_bus_out_nc_if
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_0061C_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_0061C_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:7:15
								localparam UUID_WIDTH = 1;
								// Trace: src/VX_mem_bus_if.sv:9:5
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:13:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:21:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:30:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:31:5
								// Trace: src/VX_mem_bus_if.sv:39:5
							end
							// Trace: src/VX_cache_bypass.sv:106:5
							genvar _gv_i_181;
							for (_gv_i_181 = 0; _gv_i_181 < MEM_PORTS; _gv_i_181 = _gv_i_181 + 1) begin : g_mem_bus_out_nc
								localparam i = _gv_i_181;
								// Trace: src/VX_cache_bypass.sv:107:9
								wire core_req_nc_arb_rw;
								// Trace: src/VX_cache_bypass.sv:108:9
								wire [63:0] core_req_nc_arb_byteen;
								// Trace: src/VX_cache_bypass.sv:109:9
								wire [25:0] core_req_nc_arb_addr;
								// Trace: src/VX_cache_bypass.sv:110:9
								wire [2:0] core_req_nc_arb_flags;
								// Trace: src/VX_cache_bypass.sv:111:9
								wire [511:0] core_req_nc_arb_data;
								// Trace: src/VX_cache_bypass.sv:112:9
								wire [6:0] core_req_nc_arb_tag;
								// Trace: src/VX_cache_bypass.sv:113:9
								assign {core_req_nc_arb_rw, core_req_nc_arb_addr, core_req_nc_arb_data, core_req_nc_arb_byteen, core_req_nc_arb_flags, core_req_nc_arb_tag} = core_bus_nc_arb_if[i].req_data;
								// Trace: src/VX_cache_bypass.sv:121:9
								wire [25:0] core_req_nc_arb_addr_w;
								// Trace: src/VX_cache_bypass.sv:122:9
								wire [63:0] core_req_nc_arb_byteen_w;
								// Trace: src/VX_cache_bypass.sv:123:9
								wire [511:0] core_req_nc_arb_data_w;
								// Trace: src/VX_cache_bypass.sv:124:9
								wire [511:0] core_rsp_nc_arb_data_w;
								// Trace: src/VX_cache_bypass.sv:125:9
								wire [6:0] core_req_nc_arb_tag_w;
								// Trace: src/VX_cache_bypass.sv:126:9
								wire [6:0] core_rsp_nc_arb_tag_w;
								if (1) begin : g_single_word_line
									// Trace: src/VX_cache_bypass.sv:157:13
									assign core_req_nc_arb_addr_w = core_req_nc_arb_addr;
									// Trace: src/VX_cache_bypass.sv:158:13
									assign core_req_nc_arb_byteen_w = core_req_nc_arb_byteen;
									// Trace: src/VX_cache_bypass.sv:159:13
									assign core_req_nc_arb_data_w = core_req_nc_arb_data;
									// Trace: src/VX_cache_bypass.sv:160:13
									assign core_req_nc_arb_tag_w = core_req_nc_arb_tag;
									// Trace: src/VX_cache_bypass.sv:161:13
									assign core_rsp_nc_arb_data_w = mem_bus_out_nc_if[i].rsp_data[518-:512];
									// Trace: src/VX_cache_bypass.sv:162:13
									assign core_rsp_nc_arb_tag_w = sv2v_cast_7(mem_bus_out_nc_if[i].rsp_data[6-:7]);
								end
								// Trace: src/VX_cache_bypass.sv:164:9
								assign mem_bus_out_nc_if[i].req_valid = core_bus_nc_arb_if[i].req_valid;
								// Trace: src/VX_cache_bypass.sv:165:9
								assign mem_bus_out_nc_if[i].req_data = {core_req_nc_arb_rw, core_req_nc_arb_addr_w, core_req_nc_arb_data_w, core_req_nc_arb_byteen_w, core_req_nc_arb_flags, core_req_nc_arb_tag_w};
								// Trace: src/VX_cache_bypass.sv:173:9
								assign core_bus_nc_arb_if[i].req_ready = mem_bus_out_nc_if[i].req_ready;
								// Trace: src/VX_cache_bypass.sv:174:9
								assign core_bus_nc_arb_if[i].rsp_valid = mem_bus_out_nc_if[i].rsp_valid;
								// Trace: src/VX_cache_bypass.sv:175:9
								assign core_bus_nc_arb_if[i].rsp_data = {core_rsp_nc_arb_data_w, core_rsp_nc_arb_tag_w};
								// Trace: src/VX_cache_bypass.sv:179:9
								assign mem_bus_out_nc_if[i].rsp_ready = core_bus_nc_arb_if[i].rsp_ready;
							end
							// Trace: src/VX_cache_bypass.sv:181:5
							// expanded interface instance: mem_bus_out_src_if
							localparam _param_913F6_DATA_SIZE = LINE_SIZE;
							localparam _param_913F6_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
							genvar _arr_913F6;
							for (_arr_913F6 = 0; _arr_913F6 <= (((CACHE_ENABLE ? 2 : 1) * MEM_PORTS) - 1); _arr_913F6 = _arr_913F6 + 1) begin : mem_bus_out_src_if
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_913F6_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_913F6_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:7:15
								localparam UUID_WIDTH = 1;
								// Trace: src/VX_mem_bus_if.sv:9:5
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:13:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:21:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:30:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:31:5
								// Trace: src/VX_mem_bus_if.sv:39:5
							end
							// Trace: src/VX_cache_bypass.sv:185:5
							genvar _gv_i_182;
							for (_gv_i_182 = 0; _gv_i_182 < MEM_PORTS; _gv_i_182 = _gv_i_182 + 1) begin : g_mem_bus_out_src
								localparam i = _gv_i_182;
								// Trace: src/VX_cache_bypass.sv:186:5
								assign mem_bus_out_src_if[0 + i].req_valid = mem_bus_out_nc_if[i].req_valid;
								// Trace: src/VX_cache_bypass.sv:187:5
								assign mem_bus_out_src_if[0 + i].req_data[612] = mem_bus_out_nc_if[i].req_data[612];
								// Trace: src/VX_cache_bypass.sv:188:5
								assign mem_bus_out_src_if[0 + i].req_data[611-:26] = mem_bus_out_nc_if[i].req_data[611-:26];
								// Trace: src/VX_cache_bypass.sv:189:5
								assign mem_bus_out_src_if[0 + i].req_data[585-:512] = mem_bus_out_nc_if[i].req_data[585-:512];
								// Trace: src/VX_cache_bypass.sv:190:5
								assign mem_bus_out_src_if[0 + i].req_data[73-:64] = mem_bus_out_nc_if[i].req_data[73-:64];
								// Trace: src/VX_cache_bypass.sv:191:5
								assign mem_bus_out_src_if[0 + i].req_data[9-:3] = mem_bus_out_nc_if[i].req_data[9-:3];
								if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk1
									if (1) begin : genblk1
										if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
											// Trace: src/VX_cache_bypass.sv:196:17
											assign mem_bus_out_src_if[0 + i].req_data[6-:7] = {mem_bus_out_nc_if[i].req_data[6-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_NC2_WIDTH {1'b0}}, mem_bus_out_nc_if[i].req_data[5-:6]};
										end
										else begin : genblk1
											// Trace: src/VX_cache_bypass.sv:198:17
											assign mem_bus_out_src_if[0 + i].req_data[6-:7] = {mem_bus_out_nc_if[i].req_data[6-:1], mem_bus_out_nc_if[i].req_data[(MEM_TAG_OUT_WIDTH - UUID_WIDTH) - 1:0]};
										end
									end
								end
								else begin : genblk1
									// Trace: src/VX_cache_bypass.sv:208:9
									assign mem_bus_out_src_if[0 + i].req_data[6-:7] = mem_bus_out_nc_if[i].req_data[6-:7];
								end
								// Trace: src/VX_cache_bypass.sv:211:5
								assign mem_bus_out_nc_if[i].req_ready = mem_bus_out_src_if[0 + i].req_ready;
								// Trace: src/VX_cache_bypass.sv:212:5
								assign mem_bus_out_nc_if[i].rsp_valid = mem_bus_out_src_if[0 + i].rsp_valid;
								// Trace: src/VX_cache_bypass.sv:213:5
								assign mem_bus_out_nc_if[i].rsp_data[518-:512] = mem_bus_out_src_if[0 + i].rsp_data[518-:512];
								if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk2
									if (1) begin : genblk1
										if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
											// Trace: src/VX_cache_bypass.sv:218:17
											assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[6-:1], mem_bus_out_src_if[0 + i].rsp_data[5:0]};
										end
										else begin : genblk1
											// Trace: src/VX_cache_bypass.sv:220:17
											assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[6-:1], {MEM_TAG_NC2_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[0 + i].rsp_data[5-:6]};
										end
									end
								end
								else begin : genblk2
									// Trace: src/VX_cache_bypass.sv:230:9
									assign mem_bus_out_nc_if[i].rsp_data[6-:7] = mem_bus_out_src_if[0 + i].rsp_data[6-:7];
								end
								// Trace: src/VX_cache_bypass.sv:233:5
								assign mem_bus_out_src_if[0 + i].rsp_ready = mem_bus_out_nc_if[i].rsp_ready;
								if (CACHE_ENABLE) begin : g_cache
									// Trace: src/VX_cache_bypass.sv:235:5
									assign mem_bus_out_src_if[1 + i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_valid;
									// Trace: src/VX_cache_bypass.sv:236:5
									assign mem_bus_out_src_if[1 + i].req_data[612] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[610];
									// Trace: src/VX_cache_bypass.sv:237:5
									assign mem_bus_out_src_if[1 + i].req_data[611-:26] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[609-:26];
									// Trace: src/VX_cache_bypass.sv:238:5
									assign mem_bus_out_src_if[1 + i].req_data[585-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[583-:512];
									// Trace: src/VX_cache_bypass.sv:239:5
									assign mem_bus_out_src_if[1 + i].req_data[73-:64] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[71-:64];
									// Trace: src/VX_cache_bypass.sv:240:5
									assign mem_bus_out_src_if[1 + i].req_data[9-:3] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[7-:3];
									if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk1
										if (1) begin : genblk1
											if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
												// Trace: src/VX_cache_bypass.sv:245:17
												assign mem_bus_out_src_if[1 + i].req_data[6-:7] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_IN_WIDTH {1'b0}}, Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[3-:4]};
											end
											else begin : genblk1
												// Trace: src/VX_cache_bypass.sv:247:17
												assign mem_bus_out_src_if[1 + i].req_data[6-:7] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[(MEM_TAG_OUT_WIDTH - UUID_WIDTH) - 1:0]};
											end
										end
									end
									else begin : genblk1
										// Trace: src/VX_cache_bypass.sv:257:9
										assign mem_bus_out_src_if[1 + i].req_data[6-:7] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:5];
									end
									// Trace: src/VX_cache_bypass.sv:260:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = mem_bus_out_src_if[1 + i].req_ready;
									// Trace: src/VX_cache_bypass.sv:261:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = mem_bus_out_src_if[1 + i].rsp_valid;
									// Trace: src/VX_cache_bypass.sv:262:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[516-:512] = mem_bus_out_src_if[1 + i].rsp_data[518-:512];
									if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk2
										if (1) begin : genblk1
											if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
												// Trace: src/VX_cache_bypass.sv:267:17
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[6-:1], mem_bus_out_src_if[1 + i].rsp_data[3:0]};
											end
											else begin : genblk1
												// Trace: src/VX_cache_bypass.sv:269:17
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[6-:1], {MEM_TAG_IN_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[1 + i].rsp_data[5-:6]};
											end
										end
									end
									else begin : genblk2
										// Trace: src/VX_cache_bypass.sv:279:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = mem_bus_out_src_if[1 + i].rsp_data[6-:7];
									end
									// Trace: src/VX_cache_bypass.sv:282:5
									assign mem_bus_out_src_if[1 + i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_ready;
								end
								else begin : g_no_cache
									// Trace: src/VX_cache_bypass.sv:284:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = 0;
									// Trace: src/VX_cache_bypass.sv:285:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = 0;
									// Trace: src/VX_cache_bypass.sv:286:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data = 1'sb0;
								end
							end
							// Trace: src/VX_cache_bypass.sv:289:5
							// expanded module instance: mem_bus_out_arb
							localparam _bbase_B06D0_bus_in_if = 0;
							localparam _bbase_B06D0_bus_out_if = 0;
							localparam _param_B06D0_NUM_INPUTS = (CACHE_ENABLE ? 2 : 1) * MEM_PORTS;
							localparam _param_B06D0_NUM_OUTPUTS = MEM_PORTS;
							localparam _param_B06D0_DATA_SIZE = LINE_SIZE;
							localparam _param_B06D0_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
							localparam _param_B06D0_ARBITER = "R";
							localparam _param_B06D0_REQ_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
							localparam _param_B06D0_RSP_OUT_BUF = 0;
							if (1) begin : mem_bus_out_arb
								// Trace: src/VX_mem_arb.sv:2:15
								localparam NUM_INPUTS = _param_B06D0_NUM_INPUTS;
								// Trace: src/VX_mem_arb.sv:3:15
								localparam NUM_OUTPUTS = _param_B06D0_NUM_OUTPUTS;
								// Trace: src/VX_mem_arb.sv:4:15
								localparam DATA_SIZE = _param_B06D0_DATA_SIZE;
								// Trace: src/VX_mem_arb.sv:5:15
								localparam TAG_WIDTH = _param_B06D0_TAG_WIDTH;
								// Trace: src/VX_mem_arb.sv:6:15
								localparam TAG_SEL_IDX = 0;
								// Trace: src/VX_mem_arb.sv:7:15
								localparam REQ_OUT_BUF = _param_B06D0_REQ_OUT_BUF;
								// Trace: src/VX_mem_arb.sv:8:15
								localparam RSP_OUT_BUF = _param_B06D0_RSP_OUT_BUF;
								// Trace: src/VX_mem_arb.sv:9:16
								localparam ARBITER = _param_B06D0_ARBITER;
								// Trace: src/VX_mem_arb.sv:10:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_arb.sv:11:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_arb.sv:12:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_arb.sv:14:5
								wire clk;
								// Trace: src/VX_mem_arb.sv:15:5
								wire reset;
								// Trace: src/VX_mem_arb.sv:16:5
								localparam _mbase_bus_in_if = 0;
								// Trace: src/VX_mem_arb.sv:17:5
								localparam _mbase_bus_out_if = 0;
								// Trace: src/VX_mem_arb.sv:19:5
								localparam DATA_WIDTH = 512;
								// Trace: src/VX_mem_arb.sv:20:5
								localparam LOG_NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? $clog2((NUM_INPUTS + 0) / 1) : 0);
								// Trace: src/VX_mem_arb.sv:21:5
								localparam REQ_DATAW = 606 + TAG_WIDTH;
								// Trace: src/VX_mem_arb.sv:22:5
								localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
								// Trace: src/VX_mem_arb.sv:24:5
								wire [NUM_INPUTS - 1:0] req_valid_in;
								// Trace: src/VX_mem_arb.sv:25:5
								wire [(NUM_INPUTS * REQ_DATAW) - 1:0] req_data_in;
								// Trace: src/VX_mem_arb.sv:26:5
								wire [NUM_INPUTS - 1:0] req_ready_in;
								// Trace: src/VX_mem_arb.sv:27:5
								wire [0:0] req_valid_out;
								// Trace: src/VX_mem_arb.sv:28:5
								wire [REQ_DATAW - 1:0] req_data_out;
								// Trace: src/VX_mem_arb.sv:29:5
								wire [(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1) - 1:0] req_sel_out;
								// Trace: src/VX_mem_arb.sv:30:5
								wire [0:0] req_ready_out;
								// Trace: src/VX_mem_arb.sv:31:5
								genvar _gv_i_80;
								for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
									localparam i = _gv_i_80;
									// Trace: src/VX_mem_arb.sv:32:9
									assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_valid;
									// Trace: src/VX_mem_arb.sv:33:9
									assign req_data_in[i * 613+:613] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_data;
									// Trace: src/VX_mem_arb.sv:34:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
								end
								// Trace: src/VX_mem_arb.sv:36:5
								VX_stream_arb #(
									.NUM_INPUTS(NUM_INPUTS),
									.NUM_OUTPUTS(NUM_OUTPUTS),
									.DATAW(REQ_DATAW),
									.ARBITER(ARBITER),
									.OUT_BUF(REQ_OUT_BUF)
								) req_arb(
									.clk(clk),
									.reset(reset),
									.valid_in(req_valid_in),
									.ready_in(req_ready_in),
									.data_in(req_data_in),
									.data_out(req_data_out),
									.sel_out(req_sel_out),
									.valid_out(req_valid_out),
									.ready_out(req_ready_out)
								);
								// Trace: src/VX_mem_arb.sv:53:5
								genvar _gv_i_81;
								for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
									localparam i = _gv_i_81;
									// Trace: src/VX_mem_arb.sv:54:9
									wire [TAG_WIDTH - 1:0] req_tag_out;
									// Trace: src/VX_mem_arb.sv:55:9
									VX_bits_insert #(
										.N(TAG_WIDTH),
										.S(LOG_NUM_REQS),
										.POS(TAG_SEL_IDX)
									) bits_insert(
										.data_in(req_tag_out),
										.ins_in(req_sel_out[i * 1+:1]),
										.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[6-:7])
									);
									// Trace: src/VX_mem_arb.sv:64:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
									// Trace: src/VX_mem_arb.sv:65:9
									assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[612], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[611-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[585-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[73-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[9-:3], req_tag_out} = req_data_out[i * 613+:613];
									// Trace: src/VX_mem_arb.sv:73:9
									assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
								end
								// Trace: src/VX_mem_arb.sv:75:5
								wire [NUM_INPUTS - 1:0] rsp_valid_out;
								// Trace: src/VX_mem_arb.sv:76:5
								wire [(NUM_INPUTS * RSP_DATAW) - 1:0] rsp_data_out;
								// Trace: src/VX_mem_arb.sv:77:5
								wire [NUM_INPUTS - 1:0] rsp_ready_out;
								// Trace: src/VX_mem_arb.sv:78:5
								wire [0:0] rsp_valid_in;
								// Trace: src/VX_mem_arb.sv:79:5
								wire [RSP_DATAW - 1:0] rsp_data_in;
								// Trace: src/VX_mem_arb.sv:80:5
								wire [0:0] rsp_ready_in;
								// Trace: src/VX_mem_arb.sv:81:5
								if (NUM_INPUTS > NUM_OUTPUTS) begin : g_rsp_enabled
									// Trace: src/VX_mem_arb.sv:82:9
									wire [LOG_NUM_REQS - 1:0] rsp_sel_in;
									genvar _gv_i_82;
									for (_gv_i_82 = 0; _gv_i_82 < NUM_OUTPUTS; _gv_i_82 = _gv_i_82 + 1) begin : g_rsp_data_in
										localparam i = _gv_i_82;
										// Trace: src/VX_mem_arb.sv:84:13
										wire [TAG_WIDTH - 1:0] rsp_tag_out;
										// Trace: src/VX_mem_arb.sv:85:13
										VX_bits_remove #(
											.N(TAG_WIDTH + LOG_NUM_REQS),
											.S(LOG_NUM_REQS),
											.POS(TAG_SEL_IDX)
										) bits_remove(
											.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[6-:7]),
											.sel_out(rsp_sel_in[0+:0]),
											.data_out(rsp_tag_out)
										);
										// Trace: src/VX_mem_arb.sv:94:13
										assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
										// Trace: src/VX_mem_arb.sv:95:13
										assign rsp_data_in[i * 519+:519] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[518-:512], rsp_tag_out};
										// Trace: src/VX_mem_arb.sv:96:13
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:98:9
									VX_stream_switch #(
										.NUM_INPUTS(NUM_OUTPUTS),
										.NUM_OUTPUTS(NUM_INPUTS),
										.DATAW(RSP_DATAW),
										.OUT_BUF(RSP_OUT_BUF)
									) rsp_switch(
										.clk(clk),
										.reset(reset),
										.sel_in(rsp_sel_in),
										.valid_in(rsp_valid_in),
										.ready_in(rsp_ready_in),
										.data_in(rsp_data_in),
										.data_out(rsp_data_out),
										.valid_out(rsp_valid_out),
										.ready_out(rsp_ready_out)
									);
								end
								else begin : g_passthru
									genvar _gv_i_83;
									for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
										localparam i = _gv_i_83;
										// Trace: src/VX_mem_arb.sv:116:13
										assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
										// Trace: src/VX_mem_arb.sv:117:13
										assign rsp_data_in[i * 519+:519] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
										// Trace: src/VX_mem_arb.sv:118:13
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:120:9
									VX_stream_arb #(
										.NUM_INPUTS(NUM_OUTPUTS),
										.NUM_OUTPUTS(NUM_INPUTS),
										.DATAW(RSP_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(RSP_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(rsp_valid_in),
										.ready_in(rsp_ready_in),
										.data_in(rsp_data_in),
										.data_out(rsp_data_out),
										.valid_out(rsp_valid_out),
										.ready_out(rsp_ready_out),
										.sel_out()
									);
								end
								// Trace: src/VX_mem_arb.sv:138:5
								genvar _gv_i_84;
								for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
									localparam i = _gv_i_84;
									// Trace: src/VX_mem_arb.sv:139:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
									// Trace: src/VX_mem_arb.sv:140:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
									// Trace: src/VX_mem_arb.sv:141:9
									assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_ready;
								end
							end
							assign mem_bus_out_arb.clk = clk;
							assign mem_bus_out_arb.reset = reset;
						end
						assign cache_bypass.clk = clk;
						assign cache_bypass.reset = reset;
					end
					else begin : g_no_bypass
						genvar _gv_i_167;
						for (_gv_i_167 = 0; _gv_i_167 < NUM_REQS; _gv_i_167 = _gv_i_167 + 1) begin : g_core_bus_cache_if
							localparam i = _gv_i_167;
							// Trace: src/VX_cache_wrap.sv:76:5
							assign core_bus_cache_if[i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].req_valid;
							// Trace: src/VX_cache_wrap.sv:77:5
							assign core_bus_cache_if[i].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].req_data;
							// Trace: src/VX_cache_wrap.sv:78:5
							assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].req_ready = core_bus_cache_if[i].req_ready;
							// Trace: src/VX_cache_wrap.sv:79:5
							assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].rsp_valid = core_bus_cache_if[i].rsp_valid;
							// Trace: src/VX_cache_wrap.sv:80:5
							assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].rsp_data = core_bus_cache_if[i].rsp_data;
							// Trace: src/VX_cache_wrap.sv:81:5
							assign core_bus_cache_if[i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].rsp_ready;
						end
						genvar _gv_i_168;
						for (_gv_i_168 = 0; _gv_i_168 < MEM_PORTS; _gv_i_168 = _gv_i_168 + 1) begin : g_mem_bus_tmp_if
							localparam i = _gv_i_168;
							// Trace: src/VX_cache_wrap.sv:84:5
							assign mem_bus_tmp_if[i].req_valid = mem_bus_cache_if[i].req_valid;
							// Trace: src/VX_cache_wrap.sv:85:5
							assign mem_bus_tmp_if[i].req_data = mem_bus_cache_if[i].req_data;
							// Trace: src/VX_cache_wrap.sv:86:5
							assign mem_bus_cache_if[i].req_ready = mem_bus_tmp_if[i].req_ready;
							// Trace: src/VX_cache_wrap.sv:87:5
							assign mem_bus_cache_if[i].rsp_valid = mem_bus_tmp_if[i].rsp_valid;
							// Trace: src/VX_cache_wrap.sv:88:5
							assign mem_bus_cache_if[i].rsp_data = mem_bus_tmp_if[i].rsp_data;
							// Trace: src/VX_cache_wrap.sv:89:5
							assign mem_bus_tmp_if[i].rsp_ready = mem_bus_cache_if[i].rsp_ready;
						end
					end
					// Trace: src/VX_cache_wrap.sv:92:5
					genvar _gv_i_169;
					for (_gv_i_169 = 0; _gv_i_169 < MEM_PORTS; _gv_i_169 = _gv_i_169 + 1) begin : g_mem_bus_if
						localparam i = _gv_i_169;
						if (WRITE_ENABLE) begin : g_we
							// Trace: src/VX_cache_wrap.sv:94:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
							// Trace: src/VX_cache_wrap.sv:95:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
							// Trace: src/VX_cache_wrap.sv:96:5
							assign mem_bus_tmp_if[i].req_ready = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
							// Trace: src/VX_cache_wrap.sv:97:5
							assign mem_bus_tmp_if[i].rsp_valid = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
							// Trace: src/VX_cache_wrap.sv:98:5
							assign mem_bus_tmp_if[i].rsp_data = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
							// Trace: src/VX_cache_wrap.sv:99:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
						end
						else begin : g_ro
							// Trace: src/VX_cache_wrap.sv:101:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
							// Trace: src/VX_cache_wrap.sv:102:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[612] = 0;
							// Trace: src/VX_cache_wrap.sv:103:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[611-:26] = mem_bus_tmp_if[i].req_data[611-:26];
							// Trace: src/VX_cache_wrap.sv:104:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[585-:512] = 1'sb0;
							// Trace: src/VX_cache_wrap.sv:105:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[73-:64] = 1'sb1;
							// Trace: src/VX_cache_wrap.sv:106:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[9-:3] = mem_bus_tmp_if[i].req_data[9-:3];
							// Trace: src/VX_cache_wrap.sv:107:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[6-:7] = mem_bus_tmp_if[i].req_data[6-:7];
							// Trace: src/VX_cache_wrap.sv:108:5
							assign mem_bus_tmp_if[i].req_ready = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
							// Trace: src/VX_cache_wrap.sv:109:5
							assign mem_bus_tmp_if[i].rsp_valid = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
							// Trace: src/VX_cache_wrap.sv:110:5
							assign mem_bus_tmp_if[i].rsp_data[518-:512] = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[518-:512];
							// Trace: src/VX_cache_wrap.sv:111:5
							assign mem_bus_tmp_if[i].rsp_data[6-:7] = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[6-:7];
							// Trace: src/VX_cache_wrap.sv:112:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
						end
					end
					// Trace: src/VX_cache_wrap.sv:115:5
					if (1) begin : g_passthru
						genvar _gv_i_170;
						for (_gv_i_170 = 0; _gv_i_170 < NUM_REQS; _gv_i_170 = _gv_i_170 + 1) begin : g_core_bus_cache_if
							localparam i = _gv_i_170;
							// Trace: src/VX_cache_wrap.sv:146:5
							assign core_bus_cache_if[i].req_ready = 0;
							// Trace: src/VX_cache_wrap.sv:147:5
							assign core_bus_cache_if[i].rsp_valid = 0;
							// Trace: src/VX_cache_wrap.sv:148:5
							assign core_bus_cache_if[i].rsp_data = 1'sb0;
						end
						genvar _gv_i_171;
						for (_gv_i_171 = 0; _gv_i_171 < MEM_PORTS; _gv_i_171 = _gv_i_171 + 1) begin : g_mem_bus_cache_if
							localparam i = _gv_i_171;
							// Trace: src/VX_cache_wrap.sv:151:5
							assign mem_bus_cache_if[i].req_valid = 0;
							// Trace: src/VX_cache_wrap.sv:152:5
							assign mem_bus_cache_if[i].req_data = 1'sb0;
							// Trace: src/VX_cache_wrap.sv:153:5
							assign mem_bus_cache_if[i].rsp_ready = 0;
						end
					end
				end
				assign l2cache.clk = clk;
				assign l2cache.reset = l2_reset;
				// Trace: src/VX_cluster.sv:51:5
				wire [0:0] per_socket_busy;
				// Trace: src/VX_cluster.sv:52:5
				genvar _gv_socket_id_1;
				for (_gv_socket_id_1 = 0; _gv_socket_id_1 < 1; _gv_socket_id_1 = _gv_socket_id_1 + 1) begin : g_sockets
					localparam socket_id = _gv_socket_id_1;
					// Trace: src/VX_cluster.sv:53:5
					wire [0:0] socket_reset;
					// Trace: src/VX_cluster.sv:54:5
					VX_reset_relay #(
						.N(1),
						.MAX_FANOUT(0)
					) __socket_reset(
						.clk(clk),
						.reset(reset),
						.reset_o(socket_reset)
					);
					// Trace: src/VX_cluster.sv:59:9
					// expanded interface instance: socket_dcr_bus_if
					if (1) begin : socket_dcr_bus_if
						// Trace: src/VX_dcr_bus_if.sv:2:5
						wire write_valid;
						// Trace: src/VX_dcr_bus_if.sv:3:5
						wire [11:0] write_addr;
						// Trace: src/VX_dcr_bus_if.sv:4:5
						wire [31:0] write_data;
						// Trace: src/VX_dcr_bus_if.sv:5:5
						// Trace: src/VX_dcr_bus_if.sv:10:5
					end
					// Trace: src/VX_cluster.sv:60:9
					wire is_base_dcr_addr = (Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_addr >= 12'h001) && (Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_addr < 12'h006);
					if (1) begin : genblk1
						// Trace: src/VX_cluster.sv:74:9
						assign {socket_dcr_bus_if.write_valid, socket_dcr_bus_if.write_addr, socket_dcr_bus_if.write_data} = {Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_valid && is_base_dcr_addr, Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_addr, Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_data};
					end
					// Trace: src/VX_cluster.sv:77:9
					// expanded module instance: socket
					localparam _bbase_66BD2_mem_bus_if = socket_id * VX_gpu_pkg_DCACHE_NUM_REQS;
					localparam _param_66BD2_SOCKET_ID = (CLUSTER_ID * 1) + socket_id;
					localparam _param_66BD2_INSTANCE_ID = "";
					if (1) begin : socket
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_socket.sv:2:15
						localparam SOCKET_ID = _param_66BD2_SOCKET_ID;
						// Trace: src/VX_socket.sv:3:16
						localparam INSTANCE_ID = _param_66BD2_INSTANCE_ID;
						// Trace: src/VX_socket.sv:5:5
						wire clk;
						// Trace: src/VX_socket.sv:6:5
						wire reset;
						// Trace: src/VX_socket.sv:7:5
						// removed modport instance dcr_bus_if
						// Trace: src/VX_socket.sv:8:5
						localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
						localparam VX_gpu_pkg_LSU_WORD_SIZE = 4;
						localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
						localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
						localparam _mbase_mem_bus_if = _bbase_66BD2_mem_bus_if;
						// Trace: src/VX_socket.sv:9:5
						wire busy;
						// Trace: src/VX_socket.sv:11:5
						localparam VX_gpu_pkg_ICACHE_TAG_ID_BITS = 2;
						localparam VX_gpu_pkg_ICACHE_TAG_WIDTH = 3;
						localparam VX_gpu_pkg_ICACHE_WORD_SIZE = 4;
						// expanded interface instance: per_core_icache_bus_if
						localparam _param_FD2E2_DATA_SIZE = VX_gpu_pkg_ICACHE_WORD_SIZE;
						localparam _param_FD2E2_TAG_WIDTH = VX_gpu_pkg_ICACHE_TAG_WIDTH;
						genvar _arr_FD2E2;
						for (_arr_FD2E2 = 0; _arr_FD2E2 <= 0; _arr_FD2E2 = _arr_FD2E2 + 1) begin : per_core_icache_bus_if
							// Trace: src/VX_mem_bus_if.sv:2:15
							localparam DATA_SIZE = _param_FD2E2_DATA_SIZE;
							// Trace: src/VX_mem_bus_if.sv:3:15
							localparam FLAGS_WIDTH = 3;
							// Trace: src/VX_mem_bus_if.sv:4:15
							localparam TAG_WIDTH = _param_FD2E2_TAG_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:5:15
							localparam MEM_ADDR_WIDTH = 32;
							// Trace: src/VX_mem_bus_if.sv:6:15
							localparam ADDR_WIDTH = 30;
							// Trace: src/VX_mem_bus_if.sv:7:15
							localparam UUID_WIDTH = 1;
							// Trace: src/VX_mem_bus_if.sv:9:5
							// removed localparam type tag_t
							// Trace: src/VX_mem_bus_if.sv:13:5
							// removed localparam type req_data_t
							// Trace: src/VX_mem_bus_if.sv:21:5
							// removed localparam type rsp_data_t
							// Trace: src/VX_mem_bus_if.sv:25:5
							wire req_valid;
							// Trace: src/VX_mem_bus_if.sv:26:5
							wire [72:0] req_data;
							// Trace: src/VX_mem_bus_if.sv:27:5
							wire req_ready;
							// Trace: src/VX_mem_bus_if.sv:28:5
							wire rsp_valid;
							// Trace: src/VX_mem_bus_if.sv:29:5
							wire [34:0] rsp_data;
							// Trace: src/VX_mem_bus_if.sv:30:5
							wire rsp_ready;
							// Trace: src/VX_mem_bus_if.sv:31:5
							// Trace: src/VX_mem_bus_if.sv:39:5
						end
						// Trace: src/VX_socket.sv:15:5
						localparam VX_gpu_pkg_ICACHE_LINE_SIZE = 64;
						localparam VX_gpu_pkg_ICACHE_MEM_TAG_WIDTH = 5;
						// expanded interface instance: icache_mem_bus_if
						localparam _param_063FD_DATA_SIZE = VX_gpu_pkg_ICACHE_LINE_SIZE;
						localparam _param_063FD_TAG_WIDTH = VX_gpu_pkg_ICACHE_MEM_TAG_WIDTH;
						genvar _arr_063FD;
						for (_arr_063FD = 0; _arr_063FD <= 0; _arr_063FD = _arr_063FD + 1) begin : icache_mem_bus_if
							// Trace: src/VX_mem_bus_if.sv:2:15
							localparam DATA_SIZE = _param_063FD_DATA_SIZE;
							// Trace: src/VX_mem_bus_if.sv:3:15
							localparam FLAGS_WIDTH = 3;
							// Trace: src/VX_mem_bus_if.sv:4:15
							localparam TAG_WIDTH = _param_063FD_TAG_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:5:15
							localparam MEM_ADDR_WIDTH = 32;
							// Trace: src/VX_mem_bus_if.sv:6:15
							localparam ADDR_WIDTH = 26;
							// Trace: src/VX_mem_bus_if.sv:7:15
							localparam UUID_WIDTH = 1;
							// Trace: src/VX_mem_bus_if.sv:9:5
							// removed localparam type tag_t
							// Trace: src/VX_mem_bus_if.sv:13:5
							// removed localparam type req_data_t
							// Trace: src/VX_mem_bus_if.sv:21:5
							// removed localparam type rsp_data_t
							// Trace: src/VX_mem_bus_if.sv:25:5
							wire req_valid;
							// Trace: src/VX_mem_bus_if.sv:26:5
							wire [610:0] req_data;
							// Trace: src/VX_mem_bus_if.sv:27:5
							wire req_ready;
							// Trace: src/VX_mem_bus_if.sv:28:5
							wire rsp_valid;
							// Trace: src/VX_mem_bus_if.sv:29:5
							wire [516:0] rsp_data;
							// Trace: src/VX_mem_bus_if.sv:30:5
							wire rsp_ready;
							// Trace: src/VX_mem_bus_if.sv:31:5
							// Trace: src/VX_mem_bus_if.sv:39:5
						end
						// Trace: src/VX_socket.sv:19:5
						wire [0:0] icache_reset;
						// Trace: src/VX_socket.sv:20:5
						VX_reset_relay #(
							.N(1),
							.MAX_FANOUT(0)
						) __icache_reset(
							.clk(clk),
							.reset(reset),
							.reset_o(icache_reset)
						);
						// Trace: src/VX_socket.sv:25:5
						// expanded module instance: icache
						localparam _bbase_9B047_core_bus_if = 0;
						localparam _bbase_9B047_mem_bus_if = 0;
						localparam _param_9B047_INSTANCE_ID = "";
						localparam _param_9B047_NUM_UNITS = 1;
						localparam _param_9B047_NUM_INPUTS = 1;
						localparam _param_9B047_TAG_SEL_IDX = 0;
						localparam _param_9B047_CACHE_SIZE = 16384;
						localparam _param_9B047_LINE_SIZE = VX_gpu_pkg_ICACHE_LINE_SIZE;
						localparam _param_9B047_NUM_BANKS = 1;
						localparam _param_9B047_NUM_WAYS = 4;
						localparam _param_9B047_WORD_SIZE = VX_gpu_pkg_ICACHE_WORD_SIZE;
						localparam _param_9B047_NUM_REQS = 1;
						localparam _param_9B047_MEM_PORTS = 1;
						localparam _param_9B047_CRSQ_SIZE = 2;
						localparam _param_9B047_MSHR_SIZE = 16;
						localparam _param_9B047_MRSQ_SIZE = 0;
						localparam _param_9B047_MREQ_SIZE = 4;
						localparam _param_9B047_TAG_WIDTH = VX_gpu_pkg_ICACHE_TAG_WIDTH;
						localparam _param_9B047_FLAGS_WIDTH = 0;
						localparam _param_9B047_UUID_WIDTH = 1;
						localparam _param_9B047_WRITE_ENABLE = 0;
						localparam _param_9B047_REPL_POLICY = 1;
						localparam _param_9B047_NC_ENABLE = 0;
						localparam _param_9B047_CORE_OUT_BUF = 3;
						localparam _param_9B047_MEM_OUT_BUF = 2;
						if (1) begin : icache
							// removed import VX_gpu_pkg::*;
							// Trace: src/VX_cache_cluster.sv:2:16
							localparam INSTANCE_ID = _param_9B047_INSTANCE_ID;
							// Trace: src/VX_cache_cluster.sv:3:15
							localparam NUM_UNITS = _param_9B047_NUM_UNITS;
							// Trace: src/VX_cache_cluster.sv:4:15
							localparam NUM_INPUTS = _param_9B047_NUM_INPUTS;
							// Trace: src/VX_cache_cluster.sv:5:15
							localparam TAG_SEL_IDX = _param_9B047_TAG_SEL_IDX;
							// Trace: src/VX_cache_cluster.sv:6:15
							localparam NUM_REQS = _param_9B047_NUM_REQS;
							// Trace: src/VX_cache_cluster.sv:7:15
							localparam MEM_PORTS = _param_9B047_MEM_PORTS;
							// Trace: src/VX_cache_cluster.sv:8:15
							localparam CACHE_SIZE = _param_9B047_CACHE_SIZE;
							// Trace: src/VX_cache_cluster.sv:9:15
							localparam LINE_SIZE = _param_9B047_LINE_SIZE;
							// Trace: src/VX_cache_cluster.sv:10:15
							localparam NUM_BANKS = _param_9B047_NUM_BANKS;
							// Trace: src/VX_cache_cluster.sv:11:15
							localparam NUM_WAYS = _param_9B047_NUM_WAYS;
							// Trace: src/VX_cache_cluster.sv:12:15
							localparam WORD_SIZE = _param_9B047_WORD_SIZE;
							// Trace: src/VX_cache_cluster.sv:13:15
							localparam CRSQ_SIZE = _param_9B047_CRSQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:14:15
							localparam MSHR_SIZE = _param_9B047_MSHR_SIZE;
							// Trace: src/VX_cache_cluster.sv:15:15
							localparam MRSQ_SIZE = _param_9B047_MRSQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:16:15
							localparam MREQ_SIZE = _param_9B047_MREQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:17:15
							localparam WRITE_ENABLE = _param_9B047_WRITE_ENABLE;
							// Trace: src/VX_cache_cluster.sv:18:15
							localparam WRITEBACK = 0;
							// Trace: src/VX_cache_cluster.sv:19:15
							localparam DIRTY_BYTES = 0;
							// Trace: src/VX_cache_cluster.sv:20:15
							localparam REPL_POLICY = _param_9B047_REPL_POLICY;
							// Trace: src/VX_cache_cluster.sv:21:15
							localparam UUID_WIDTH = _param_9B047_UUID_WIDTH;
							// Trace: src/VX_cache_cluster.sv:22:15
							localparam TAG_WIDTH = _param_9B047_TAG_WIDTH;
							// Trace: src/VX_cache_cluster.sv:23:15
							localparam FLAGS_WIDTH = _param_9B047_FLAGS_WIDTH;
							// Trace: src/VX_cache_cluster.sv:24:15
							localparam NC_ENABLE = _param_9B047_NC_ENABLE;
							// Trace: src/VX_cache_cluster.sv:25:15
							localparam CORE_OUT_BUF = _param_9B047_CORE_OUT_BUF;
							// Trace: src/VX_cache_cluster.sv:26:15
							localparam MEM_OUT_BUF = _param_9B047_MEM_OUT_BUF;
							// Trace: src/VX_cache_cluster.sv:28:5
							wire clk;
							// Trace: src/VX_cache_cluster.sv:29:5
							wire reset;
							// Trace: src/VX_cache_cluster.sv:30:5
							localparam _mbase_core_bus_if = 0;
							// Trace: src/VX_cache_cluster.sv:31:5
							localparam _mbase_mem_bus_if = 0;
							// Trace: src/VX_cache_cluster.sv:33:5
							localparam NUM_CACHES = NUM_UNITS;
							// Trace: src/VX_cache_cluster.sv:34:5
							localparam PASSTHRU = 1'd0;
							// Trace: src/VX_cache_cluster.sv:35:5
							localparam ARB_TAG_WIDTH = 3;
							// Trace: src/VX_cache_cluster.sv:36:5
							localparam CACHE_MEM_TAG_WIDTH = 5;
							// Trace: src/VX_cache_cluster.sv:38:5
							localparam BYPASS_TAG_WIDTH = 7;
							// Trace: src/VX_cache_cluster.sv:40:5
							localparam NC_TAG_WIDTH = 8;
							// Trace: src/VX_cache_cluster.sv:41:5
							localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
							// Trace: src/VX_cache_cluster.sv:42:5
							// expanded interface instance: cache_mem_bus_if
							localparam _param_A4879_DATA_SIZE = LINE_SIZE;
							localparam _param_A4879_TAG_WIDTH = MEM_TAG_WIDTH;
							genvar _arr_A4879;
							for (_arr_A4879 = 0; _arr_A4879 <= 0; _arr_A4879 = _arr_A4879 + 1) begin : cache_mem_bus_if
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_A4879_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_A4879_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:7:15
								localparam UUID_WIDTH = 1;
								// Trace: src/VX_mem_bus_if.sv:9:5
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:13:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:21:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire [610:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire [516:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:30:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:31:5
								// Trace: src/VX_mem_bus_if.sv:39:5
							end
							// Trace: src/VX_cache_cluster.sv:46:5
							// expanded interface instance: arb_core_bus_if
							localparam _param_F9BC9_DATA_SIZE = WORD_SIZE;
							localparam _param_F9BC9_TAG_WIDTH = ARB_TAG_WIDTH;
							genvar _arr_F9BC9;
							for (_arr_F9BC9 = 0; _arr_F9BC9 <= 0; _arr_F9BC9 = _arr_F9BC9 + 1) begin : arb_core_bus_if
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_F9BC9_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_F9BC9_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 30;
								// Trace: src/VX_mem_bus_if.sv:7:15
								localparam UUID_WIDTH = 1;
								// Trace: src/VX_mem_bus_if.sv:9:5
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:13:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:21:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire [72:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire [34:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:30:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:31:5
								// Trace: src/VX_mem_bus_if.sv:39:5
							end
							// Trace: src/VX_cache_cluster.sv:50:5
							genvar _gv_i_65;
							for (_gv_i_65 = 0; _gv_i_65 < NUM_REQS; _gv_i_65 = _gv_i_65 + 1) begin : g_core_arb
								localparam i = _gv_i_65;
								// Trace: src/VX_cache_cluster.sv:51:9
								// expanded interface instance: core_bus_tmp_if
								localparam _param_A62F7_DATA_SIZE = WORD_SIZE;
								localparam _param_A62F7_TAG_WIDTH = TAG_WIDTH;
								genvar _arr_A62F7;
								for (_arr_A62F7 = 0; _arr_A62F7 <= 0; _arr_A62F7 = _arr_A62F7 + 1) begin : core_bus_tmp_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_A62F7_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_A62F7_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 30;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [72:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [34:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								// Trace: src/VX_cache_cluster.sv:55:9
								// expanded interface instance: arb_core_bus_tmp_if
								localparam _param_E788B_DATA_SIZE = WORD_SIZE;
								localparam _param_E788B_TAG_WIDTH = ARB_TAG_WIDTH;
								genvar _arr_E788B;
								for (_arr_E788B = 0; _arr_E788B <= 0; _arr_E788B = _arr_E788B + 1) begin : arb_core_bus_tmp_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_E788B_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_E788B_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 30;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [72:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [34:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								genvar _gv_j_6;
								for (_gv_j_6 = 0; _gv_j_6 < NUM_INPUTS; _gv_j_6 = _gv_j_6 + 1) begin : g_core_bus_tmp_if
									localparam j = _gv_j_6;
									// Trace: src/VX_cache_cluster.sv:60:5
									assign core_bus_tmp_if[j].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_valid;
									// Trace: src/VX_cache_cluster.sv:61:5
									assign core_bus_tmp_if[j].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_data;
									// Trace: src/VX_cache_cluster.sv:62:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_ready = core_bus_tmp_if[j].req_ready;
									// Trace: src/VX_cache_cluster.sv:63:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_valid = core_bus_tmp_if[j].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:64:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_data = core_bus_tmp_if[j].rsp_data;
									// Trace: src/VX_cache_cluster.sv:65:5
									assign core_bus_tmp_if[j].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_ready;
								end
								// Trace: src/VX_cache_cluster.sv:67:9
								// expanded module instance: core_arb
								localparam _bbase_856A9_bus_in_if = 0;
								localparam _bbase_856A9_bus_out_if = 0;
								localparam _param_856A9_NUM_INPUTS = NUM_INPUTS;
								localparam _param_856A9_NUM_OUTPUTS = NUM_CACHES;
								localparam _param_856A9_DATA_SIZE = WORD_SIZE;
								localparam _param_856A9_TAG_WIDTH = TAG_WIDTH;
								localparam _param_856A9_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_856A9_ARBITER = "R";
								localparam _param_856A9_REQ_OUT_BUF = 0;
								localparam _param_856A9_RSP_OUT_BUF = 0;
								if (1) begin : core_arb
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_856A9_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = _param_856A9_NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_856A9_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_856A9_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_856A9_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_856A9_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_856A9_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:16
									localparam ARBITER = _param_856A9_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 30;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 0;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 73;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = 35;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [0:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [72:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [0:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [72:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_80;
									for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
										localparam i = _gv_i_80;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 73+:73] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_81;
									for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
										localparam i = _gv_i_81;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [2:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										VX_bits_insert #(
											.N(TAG_WIDTH),
											.S(LOG_NUM_REQS),
											.POS(TAG_SEL_IDX)
										) bits_insert(
											.data_in(req_tag_out),
											.ins_in(req_sel_out[i+:1]),
											.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[2-:3])
										);
										// Trace: src/VX_mem_arb.sv:64:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:65:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[72], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[71-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[41-:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[9-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[5-:3], req_tag_out} = req_data_out[i * 73+:73];
										// Trace: src/VX_mem_arb.sv:73:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
									end
									// Trace: src/VX_mem_arb.sv:75:5
									wire [0:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:76:5
									wire [34:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:77:5
									wire [0:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:78:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:79:5
									wire [34:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:81:5
									if (1) begin : g_passthru
										genvar _gv_i_83;
										for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_83;
											// Trace: src/VX_mem_arb.sv:116:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:117:13
											assign rsp_data_in[i * 35+:35] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
											// Trace: src/VX_mem_arb.sv:118:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:120:9
										VX_stream_arb #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.ARBITER(ARBITER),
											.OUT_BUF(RSP_OUT_BUF)
										) req_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
									end
									// Trace: src/VX_mem_arb.sv:138:5
									genvar _gv_i_84;
									for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
										localparam i = _gv_i_84;
										// Trace: src/VX_mem_arb.sv:139:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:140:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 35+:35];
										// Trace: src/VX_mem_arb.sv:141:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign core_arb.clk = clk;
								assign core_arb.reset = reset;
								genvar _gv_k_1;
								for (_gv_k_1 = 0; _gv_k_1 < NUM_CACHES; _gv_k_1 = _gv_k_1 + 1) begin : g_arb_core_bus_if
									localparam k = _gv_k_1;
									// Trace: src/VX_cache_cluster.sv:83:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].req_valid = arb_core_bus_tmp_if[k].req_valid;
									// Trace: src/VX_cache_cluster.sv:84:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].req_data = arb_core_bus_tmp_if[k].req_data;
									// Trace: src/VX_cache_cluster.sv:85:5
									assign arb_core_bus_tmp_if[k].req_ready = arb_core_bus_if[(k * NUM_REQS) + i].req_ready;
									// Trace: src/VX_cache_cluster.sv:86:5
									assign arb_core_bus_tmp_if[k].rsp_valid = arb_core_bus_if[(k * NUM_REQS) + i].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:87:5
									assign arb_core_bus_tmp_if[k].rsp_data = arb_core_bus_if[(k * NUM_REQS) + i].rsp_data;
									// Trace: src/VX_cache_cluster.sv:88:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].rsp_ready = arb_core_bus_tmp_if[k].rsp_ready;
								end
							end
							// Trace: src/VX_cache_cluster.sv:91:6
							genvar _gv_i_66;
							for (_gv_i_66 = 0; _gv_i_66 < NUM_CACHES; _gv_i_66 = _gv_i_66 + 1) begin : g_cache_wrap
								localparam i = _gv_i_66;
								// Trace: src/VX_cache_cluster.sv:92:9
								// expanded module instance: cache_wrap
								localparam _bbase_665FE_core_bus_if = i * NUM_REQS;
								localparam _bbase_665FE_mem_bus_if = i * MEM_PORTS;
								localparam _param_665FE_INSTANCE_ID = "";
								localparam _param_665FE_CACHE_SIZE = CACHE_SIZE;
								localparam _param_665FE_LINE_SIZE = LINE_SIZE;
								localparam _param_665FE_NUM_BANKS = NUM_BANKS;
								localparam _param_665FE_NUM_WAYS = NUM_WAYS;
								localparam _param_665FE_WORD_SIZE = WORD_SIZE;
								localparam _param_665FE_NUM_REQS = NUM_REQS;
								localparam _param_665FE_MEM_PORTS = MEM_PORTS;
								localparam _param_665FE_WRITE_ENABLE = WRITE_ENABLE;
								localparam _param_665FE_WRITEBACK = WRITEBACK;
								localparam _param_665FE_DIRTY_BYTES = DIRTY_BYTES;
								localparam _param_665FE_REPL_POLICY = REPL_POLICY;
								localparam _param_665FE_CRSQ_SIZE = CRSQ_SIZE;
								localparam _param_665FE_MSHR_SIZE = MSHR_SIZE;
								localparam _param_665FE_MRSQ_SIZE = MRSQ_SIZE;
								localparam _param_665FE_MREQ_SIZE = MREQ_SIZE;
								localparam _param_665FE_UUID_WIDTH = UUID_WIDTH;
								localparam _param_665FE_TAG_WIDTH = ARB_TAG_WIDTH;
								localparam _param_665FE_FLAGS_WIDTH = FLAGS_WIDTH;
								localparam _param_665FE_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_665FE_CORE_OUT_BUF = CORE_OUT_BUF;
								localparam _param_665FE_MEM_OUT_BUF = MEM_OUT_BUF;
								localparam _param_665FE_NC_ENABLE = NC_ENABLE;
								localparam _param_665FE_PASSTHRU = PASSTHRU;
								if (1) begin : cache_wrap
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_cache_wrap.sv:2:16
									localparam INSTANCE_ID = _param_665FE_INSTANCE_ID;
									// Trace: src/VX_cache_wrap.sv:3:15
									localparam TAG_SEL_IDX = _param_665FE_TAG_SEL_IDX;
									// Trace: src/VX_cache_wrap.sv:4:15
									localparam NUM_REQS = _param_665FE_NUM_REQS;
									// Trace: src/VX_cache_wrap.sv:5:15
									localparam MEM_PORTS = _param_665FE_MEM_PORTS;
									// Trace: src/VX_cache_wrap.sv:6:15
									localparam CACHE_SIZE = _param_665FE_CACHE_SIZE;
									// Trace: src/VX_cache_wrap.sv:7:15
									localparam LINE_SIZE = _param_665FE_LINE_SIZE;
									// Trace: src/VX_cache_wrap.sv:8:15
									localparam NUM_BANKS = _param_665FE_NUM_BANKS;
									// Trace: src/VX_cache_wrap.sv:9:15
									localparam NUM_WAYS = _param_665FE_NUM_WAYS;
									// Trace: src/VX_cache_wrap.sv:10:15
									localparam WORD_SIZE = _param_665FE_WORD_SIZE;
									// Trace: src/VX_cache_wrap.sv:11:15
									localparam CRSQ_SIZE = _param_665FE_CRSQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:12:15
									localparam MSHR_SIZE = _param_665FE_MSHR_SIZE;
									// Trace: src/VX_cache_wrap.sv:13:15
									localparam MRSQ_SIZE = _param_665FE_MRSQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:14:15
									localparam MREQ_SIZE = _param_665FE_MREQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:15:15
									localparam WRITE_ENABLE = _param_665FE_WRITE_ENABLE;
									// Trace: src/VX_cache_wrap.sv:16:15
									localparam WRITEBACK = _param_665FE_WRITEBACK;
									// Trace: src/VX_cache_wrap.sv:17:15
									localparam DIRTY_BYTES = _param_665FE_DIRTY_BYTES;
									// Trace: src/VX_cache_wrap.sv:18:15
									localparam REPL_POLICY = _param_665FE_REPL_POLICY;
									// Trace: src/VX_cache_wrap.sv:19:15
									localparam UUID_WIDTH = _param_665FE_UUID_WIDTH;
									// Trace: src/VX_cache_wrap.sv:20:15
									localparam TAG_WIDTH = _param_665FE_TAG_WIDTH;
									// Trace: src/VX_cache_wrap.sv:21:15
									localparam FLAGS_WIDTH = _param_665FE_FLAGS_WIDTH;
									// Trace: src/VX_cache_wrap.sv:22:15
									localparam NC_ENABLE = _param_665FE_NC_ENABLE;
									// Trace: src/VX_cache_wrap.sv:23:15
									localparam PASSTHRU = _param_665FE_PASSTHRU;
									// Trace: src/VX_cache_wrap.sv:24:15
									localparam CORE_OUT_BUF = _param_665FE_CORE_OUT_BUF;
									// Trace: src/VX_cache_wrap.sv:25:15
									localparam MEM_OUT_BUF = _param_665FE_MEM_OUT_BUF;
									// Trace: src/VX_cache_wrap.sv:27:5
									wire clk;
									// Trace: src/VX_cache_wrap.sv:28:5
									wire reset;
									// Trace: src/VX_cache_wrap.sv:29:5
									localparam _mbase_core_bus_if = _bbase_665FE_core_bus_if;
									// Trace: src/VX_cache_wrap.sv:30:5
									localparam _mbase_mem_bus_if = _bbase_665FE_mem_bus_if;
									// Trace: src/VX_cache_wrap.sv:32:5
									localparam CACHE_MEM_TAG_WIDTH = 5;
									// Trace: src/VX_cache_wrap.sv:34:5
									localparam BYPASS_TAG_WIDTH = 7;
									// Trace: src/VX_cache_wrap.sv:36:5
									localparam NC_TAG_WIDTH = 8;
									// Trace: src/VX_cache_wrap.sv:37:5
									localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
									// Trace: src/VX_cache_wrap.sv:38:5
									localparam BYPASS_ENABLE = 1'd0;
									// Trace: src/VX_cache_wrap.sv:39:5
									// expanded interface instance: core_bus_cache_if
									localparam _param_24C1C_DATA_SIZE = WORD_SIZE;
									localparam _param_24C1C_TAG_WIDTH = TAG_WIDTH;
									genvar _arr_24C1C;
									for (_arr_24C1C = 0; _arr_24C1C <= 0; _arr_24C1C = _arr_24C1C + 1) begin : core_bus_cache_if
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_24C1C_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_24C1C_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_mem_bus_if.sv:7:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_mem_bus_if.sv:9:5
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:21:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire [72:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire [34:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:30:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:31:5
										// Trace: src/VX_mem_bus_if.sv:39:5
									end
									// Trace: src/VX_cache_wrap.sv:43:5
									// expanded interface instance: mem_bus_cache_if
									localparam _param_D895D_DATA_SIZE = LINE_SIZE;
									localparam _param_D895D_TAG_WIDTH = CACHE_MEM_TAG_WIDTH;
									genvar _arr_D895D;
									for (_arr_D895D = 0; _arr_D895D <= 0; _arr_D895D = _arr_D895D + 1) begin : mem_bus_cache_if
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_D895D_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_D895D_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 26;
										// Trace: src/VX_mem_bus_if.sv:7:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_mem_bus_if.sv:9:5
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:21:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire [610:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire [516:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:30:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:31:5
										// Trace: src/VX_mem_bus_if.sv:39:5
									end
									// Trace: src/VX_cache_wrap.sv:47:5
									// expanded interface instance: mem_bus_tmp_if
									localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
									localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
									genvar _arr_4FE36;
									for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 26;
										// Trace: src/VX_mem_bus_if.sv:7:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_mem_bus_if.sv:9:5
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:21:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire [610:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire [516:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:30:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:31:5
										// Trace: src/VX_mem_bus_if.sv:39:5
									end
									// Trace: src/VX_cache_wrap.sv:51:5
									if (BYPASS_ENABLE) begin : g_bypass
										// Trace: src/VX_cache_wrap.sv:52:9
										// expanded module instance: cache_bypass
										localparam _bbase_714AA_core_bus_in_if = i * NUM_REQS;
										localparam _bbase_714AA_core_bus_out_if = 0;
										localparam _bbase_714AA_mem_bus_in_if = 0;
										localparam _bbase_714AA_mem_bus_out_if = 0;
										localparam _param_714AA_NUM_REQS = NUM_REQS;
										localparam _param_714AA_MEM_PORTS = MEM_PORTS;
										localparam _param_714AA_TAG_SEL_IDX = TAG_SEL_IDX;
										localparam _param_714AA_CACHE_ENABLE = !PASSTHRU;
										localparam _param_714AA_WORD_SIZE = WORD_SIZE;
										localparam _param_714AA_LINE_SIZE = LINE_SIZE;
										localparam _param_714AA_CORE_ADDR_WIDTH = 30;
										localparam _param_714AA_CORE_TAG_WIDTH = TAG_WIDTH;
										localparam _param_714AA_MEM_ADDR_WIDTH = 26;
										localparam _param_714AA_MEM_TAG_IN_WIDTH = CACHE_MEM_TAG_WIDTH;
										localparam _param_714AA_UUID_WIDTH = UUID_WIDTH;
										localparam _param_714AA_CORE_OUT_BUF = CORE_OUT_BUF;
										localparam _param_714AA_MEM_OUT_BUF = MEM_OUT_BUF;
										if (1) begin : cache_bypass
											// Trace: src/VX_cache_bypass.sv:2:15
											localparam NUM_REQS = _param_714AA_NUM_REQS;
											// Trace: src/VX_cache_bypass.sv:3:15
											localparam MEM_PORTS = _param_714AA_MEM_PORTS;
											// Trace: src/VX_cache_bypass.sv:4:15
											localparam TAG_SEL_IDX = _param_714AA_TAG_SEL_IDX;
											// Trace: src/VX_cache_bypass.sv:5:15
											localparam CACHE_ENABLE = _param_714AA_CACHE_ENABLE;
											// Trace: src/VX_cache_bypass.sv:6:15
											localparam WORD_SIZE = _param_714AA_WORD_SIZE;
											// Trace: src/VX_cache_bypass.sv:7:15
											localparam LINE_SIZE = _param_714AA_LINE_SIZE;
											// Trace: src/VX_cache_bypass.sv:8:15
											localparam CORE_ADDR_WIDTH = _param_714AA_CORE_ADDR_WIDTH;
											// Trace: src/VX_cache_bypass.sv:9:15
											localparam CORE_TAG_WIDTH = _param_714AA_CORE_TAG_WIDTH;
											// Trace: src/VX_cache_bypass.sv:10:15
											localparam MEM_ADDR_WIDTH = _param_714AA_MEM_ADDR_WIDTH;
											// Trace: src/VX_cache_bypass.sv:11:15
											localparam MEM_TAG_IN_WIDTH = _param_714AA_MEM_TAG_IN_WIDTH;
											// Trace: src/VX_cache_bypass.sv:12:15
											localparam UUID_WIDTH = _param_714AA_UUID_WIDTH;
											// Trace: src/VX_cache_bypass.sv:13:15
											localparam CORE_OUT_BUF = _param_714AA_CORE_OUT_BUF;
											// Trace: src/VX_cache_bypass.sv:14:15
											localparam MEM_OUT_BUF = _param_714AA_MEM_OUT_BUF;
											// Trace: src/VX_cache_bypass.sv:16:5
											wire clk;
											// Trace: src/VX_cache_bypass.sv:17:5
											wire reset;
											// Trace: src/VX_cache_bypass.sv:18:5
											localparam _mbase_core_bus_in_if = _bbase_714AA_core_bus_in_if;
											// Trace: src/VX_cache_bypass.sv:19:5
											localparam _mbase_core_bus_out_if = 0;
											// Trace: src/VX_cache_bypass.sv:20:5
											localparam _mbase_mem_bus_in_if = 0;
											// Trace: src/VX_cache_bypass.sv:21:5
											localparam _mbase_mem_bus_out_if = 0;
											// Trace: src/VX_cache_bypass.sv:23:5
											localparam DIRECT_PASSTHRU = (!CACHE_ENABLE && 1'd0) && 1'd1;
											// Trace: src/VX_cache_bypass.sv:24:5
											localparam CORE_DATA_WIDTH = 32;
											// Trace: src/VX_cache_bypass.sv:25:5
											localparam WORDS_PER_LINE = 16;
											// Trace: src/VX_cache_bypass.sv:26:5
											localparam WSEL_BITS = 4;
											// Trace: src/VX_cache_bypass.sv:27:5
											localparam CORE_TAG_ID_WIDTH = 2;
											// Trace: src/VX_cache_bypass.sv:28:5
											localparam MEM_TAG_ID_WIDTH = 2;
											// Trace: src/VX_cache_bypass.sv:29:5
											localparam MEM_TAG_NC1_WIDTH = 3;
											// Trace: src/VX_cache_bypass.sv:30:5
											localparam MEM_TAG_NC2_WIDTH = 7;
											// Trace: src/VX_cache_bypass.sv:31:5
											localparam MEM_TAG_OUT_WIDTH = (CACHE_ENABLE ? MEM_TAG_NC2_WIDTH : MEM_TAG_NC2_WIDTH);
											// Trace: src/VX_cache_bypass.sv:32:5
											// expanded interface instance: core_bus_nc_switch_if
											localparam _param_95306_DATA_SIZE = WORD_SIZE;
											localparam _param_95306_TAG_WIDTH = CORE_TAG_WIDTH;
											genvar _arr_95306;
											for (_arr_95306 = 0; _arr_95306 <= (((CACHE_ENABLE ? 2 : 1) * NUM_REQS) - 1); _arr_95306 = _arr_95306 + 1) begin : core_bus_nc_switch_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_95306_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_95306_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [72:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [34:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:36:5
											wire [0:0] core_req_nc_sel;
											// Trace: src/VX_cache_bypass.sv:37:5
											genvar _gv_i_179;
											for (_gv_i_179 = 0; _gv_i_179 < NUM_REQS; _gv_i_179 = _gv_i_179 + 1) begin : g_core_req_is_nc
												localparam i = _gv_i_179;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:39:13
													assign core_req_nc_sel[i] = ~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_in_if].req_data[4];
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:41:13
													assign core_req_nc_sel[i] = 1'b0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:44:5
											// expanded module instance: core_bus_nc_switch
											localparam _bbase_69FDB_bus_in_if = i * NUM_REQS;
											localparam _bbase_69FDB_bus_out_if = 0;
											localparam _param_69FDB_NUM_INPUTS = NUM_REQS;
											localparam _param_69FDB_NUM_OUTPUTS = (CACHE_ENABLE ? 2 : 1) * NUM_REQS;
											localparam _param_69FDB_DATA_SIZE = WORD_SIZE;
											localparam _param_69FDB_TAG_WIDTH = CORE_TAG_WIDTH;
											localparam _param_69FDB_ARBITER = "R";
											localparam _param_69FDB_REQ_OUT_BUF = 0;
											localparam _param_69FDB_RSP_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
											if (1) begin : core_bus_nc_switch
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_switch.sv:2:15
												localparam NUM_INPUTS = _param_69FDB_NUM_INPUTS;
												// Trace: src/VX_mem_switch.sv:3:15
												localparam NUM_OUTPUTS = _param_69FDB_NUM_OUTPUTS;
												// Trace: src/VX_mem_switch.sv:4:15
												localparam DATA_SIZE = _param_69FDB_DATA_SIZE;
												// Trace: src/VX_mem_switch.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_switch.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_switch.sv:7:15
												localparam TAG_WIDTH = _param_69FDB_TAG_WIDTH;
												// Trace: src/VX_mem_switch.sv:8:15
												localparam REQ_OUT_BUF = _param_69FDB_REQ_OUT_BUF;
												// Trace: src/VX_mem_switch.sv:9:15
												localparam RSP_OUT_BUF = _param_69FDB_RSP_OUT_BUF;
												// Trace: src/VX_mem_switch.sv:10:16
												localparam ARBITER = _param_69FDB_ARBITER;
												// Trace: src/VX_mem_switch.sv:11:15
												localparam NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
												// Trace: src/VX_mem_switch.sv:12:15
												localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
												// Trace: src/VX_mem_switch.sv:13:15
												localparam LOG_NUM_REQS = $clog2(NUM_REQS);
												// Trace: src/VX_mem_switch.sv:15:5
												wire clk;
												// Trace: src/VX_mem_switch.sv:16:5
												wire reset;
												// Trace: src/VX_mem_switch.sv:17:5
												wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] bus_sel;
												// Trace: src/VX_mem_switch.sv:18:5
												localparam _mbase_bus_in_if = _bbase_69FDB_bus_in_if;
												// Trace: src/VX_mem_switch.sv:19:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_switch.sv:21:5
												localparam DATA_WIDTH = 32;
												// Trace: src/VX_mem_switch.sv:22:5
												localparam REQ_DATAW = 73;
												// Trace: src/VX_mem_switch.sv:23:5
												localparam RSP_DATAW = 35;
												// Trace: src/VX_mem_switch.sv:24:5
												wire [0:0] req_valid_in;
												// Trace: src/VX_mem_switch.sv:25:5
												wire [72:0] req_data_in;
												// Trace: src/VX_mem_switch.sv:26:5
												wire [0:0] req_ready_in;
												// Trace: src/VX_mem_switch.sv:27:5
												wire [NUM_OUTPUTS - 1:0] req_valid_out;
												// Trace: src/VX_mem_switch.sv:28:5
												wire [(NUM_OUTPUTS * 73) - 1:0] req_data_out;
												// Trace: src/VX_mem_switch.sv:29:5
												wire [NUM_OUTPUTS - 1:0] req_ready_out;
												// Trace: src/VX_mem_switch.sv:30:5
												genvar _gv_i_154;
												for (_gv_i_154 = 0; _gv_i_154 < NUM_INPUTS; _gv_i_154 = _gv_i_154 + 1) begin : g_req_data_in
													localparam i = _gv_i_154;
													// Trace: src/VX_mem_switch.sv:31:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_switch.sv:32:9
													assign req_data_in[i * 73+:73] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_switch.sv:33:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_switch.sv:35:5
												VX_stream_switch #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.OUT_BUF(REQ_OUT_BUF)
												) req_switch(
													.clk(clk),
													.reset(reset),
													.sel_in(bus_sel),
													.valid_in(req_valid_in),
													.data_in(req_data_in),
													.ready_in(req_ready_in),
													.valid_out(req_valid_out),
													.data_out(req_data_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_switch.sv:51:5
												genvar _gv_i_155;
												for (_gv_i_155 = 0; _gv_i_155 < NUM_OUTPUTS; _gv_i_155 = _gv_i_155 + 1) begin : g_req_data_out
													localparam i = _gv_i_155;
													// Trace: src/VX_mem_switch.sv:52:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_switch.sv:53:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_data = req_data_out[i * 73+:73];
													// Trace: src/VX_mem_switch.sv:54:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_ready;
												end
												// Trace: src/VX_mem_switch.sv:56:5
												wire [NUM_OUTPUTS - 1:0] rsp_valid_in;
												// Trace: src/VX_mem_switch.sv:57:5
												wire [(NUM_OUTPUTS * 35) - 1:0] rsp_data_in;
												// Trace: src/VX_mem_switch.sv:58:5
												wire [NUM_OUTPUTS - 1:0] rsp_ready_in;
												// Trace: src/VX_mem_switch.sv:59:5
												wire [0:0] rsp_valid_out;
												// Trace: src/VX_mem_switch.sv:60:5
												wire [34:0] rsp_data_out;
												// Trace: src/VX_mem_switch.sv:61:5
												wire [0:0] rsp_ready_out;
												// Trace: src/VX_mem_switch.sv:62:5
												genvar _gv_i_156;
												for (_gv_i_156 = 0; _gv_i_156 < NUM_OUTPUTS; _gv_i_156 = _gv_i_156 + 1) begin : g_rsp_data_in
													localparam i = _gv_i_156;
													// Trace: src/VX_mem_switch.sv:63:9
													assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_valid;
													// Trace: src/VX_mem_switch.sv:64:9
													assign rsp_data_in[i * 35+:35] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_data;
													// Trace: src/VX_mem_switch.sv:65:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
												end
												// Trace: src/VX_mem_switch.sv:67:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_OUTPUTS),
													.NUM_OUTPUTS(NUM_INPUTS),
													.DATAW(RSP_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(RSP_OUT_BUF)
												) rsp_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(rsp_valid_in),
													.data_in(rsp_data_in),
													.ready_in(rsp_ready_in),
													.valid_out(rsp_valid_out),
													.data_out(rsp_data_out),
													.ready_out(rsp_ready_out),
													.sel_out()
												);
												// Trace: src/VX_mem_switch.sv:84:5
												genvar _gv_i_157;
												for (_gv_i_157 = 0; _gv_i_157 < NUM_INPUTS; _gv_i_157 = _gv_i_157 + 1) begin : g_rsp_data_out
													localparam i = _gv_i_157;
													// Trace: src/VX_mem_switch.sv:85:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_switch.sv:86:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 35+:35];
													// Trace: src/VX_mem_switch.sv:87:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign core_bus_nc_switch.clk = clk;
											assign core_bus_nc_switch.reset = reset;
											assign core_bus_nc_switch.bus_sel = core_req_nc_sel;
											// Trace: src/VX_cache_bypass.sv:59:5
											// expanded interface instance: core_bus_in_nc_if
											localparam _param_C0263_DATA_SIZE = WORD_SIZE;
											localparam _param_C0263_TAG_WIDTH = CORE_TAG_WIDTH;
											genvar _arr_C0263;
											for (_arr_C0263 = 0; _arr_C0263 <= 0; _arr_C0263 = _arr_C0263 + 1) begin : core_bus_in_nc_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_C0263_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_C0263_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [72:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [34:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:63:5
											genvar _gv_i_180;
											for (_gv_i_180 = 0; _gv_i_180 < NUM_REQS; _gv_i_180 = _gv_i_180 + 1) begin : g_core_bus_nc_switch_if
												localparam i = _gv_i_180;
												// Trace: src/VX_cache_bypass.sv:64:9
												assign core_bus_in_nc_if[i].req_valid = core_bus_nc_switch_if[0 + i].req_valid;
												// Trace: src/VX_cache_bypass.sv:65:9
												assign core_bus_in_nc_if[i].req_data = core_bus_nc_switch_if[0 + i].req_data;
												// Trace: src/VX_cache_bypass.sv:66:9
												assign core_bus_nc_switch_if[0 + i].req_ready = core_bus_in_nc_if[i].req_ready;
												// Trace: src/VX_cache_bypass.sv:67:9
												assign core_bus_nc_switch_if[0 + i].rsp_valid = core_bus_in_nc_if[i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:68:9
												assign core_bus_nc_switch_if[0 + i].rsp_data = core_bus_in_nc_if[i].rsp_data;
												// Trace: src/VX_cache_bypass.sv:69:9
												assign core_bus_in_nc_if[i].rsp_ready = core_bus_nc_switch_if[0 + i].rsp_ready;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:71:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = core_bus_nc_switch_if[1 + i].req_valid;
													// Trace: src/VX_cache_bypass.sv:72:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = core_bus_nc_switch_if[1 + i].req_data;
													// Trace: src/VX_cache_bypass.sv:73:13
													assign core_bus_nc_switch_if[1 + i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_ready;
													// Trace: src/VX_cache_bypass.sv:74:13
													assign core_bus_nc_switch_if[1 + i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_valid;
													// Trace: src/VX_cache_bypass.sv:75:13
													assign core_bus_nc_switch_if[1 + i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_data;
													// Trace: src/VX_cache_bypass.sv:76:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = core_bus_nc_switch_if[1 + i].rsp_ready;
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:78:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = 0;
													// Trace: src/VX_cache_bypass.sv:79:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = 1'sb0;
													// Trace: src/VX_cache_bypass.sv:80:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = 0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:83:5
											// expanded interface instance: core_bus_nc_arb_if
											localparam _param_D50AC_DATA_SIZE = WORD_SIZE;
											localparam _param_D50AC_TAG_WIDTH = MEM_TAG_NC1_WIDTH;
											genvar _arr_D50AC;
											for (_arr_D50AC = 0; _arr_D50AC <= 0; _arr_D50AC = _arr_D50AC + 1) begin : core_bus_nc_arb_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_D50AC_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_D50AC_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [72:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [34:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:87:5
											// expanded module instance: core_bus_nc_arb
											localparam _bbase_1376F_bus_in_if = 0;
											localparam _bbase_1376F_bus_out_if = 0;
											localparam _param_1376F_NUM_INPUTS = NUM_REQS;
											localparam _param_1376F_NUM_OUTPUTS = MEM_PORTS;
											localparam _param_1376F_DATA_SIZE = WORD_SIZE;
											localparam _param_1376F_TAG_WIDTH = CORE_TAG_WIDTH;
											localparam _param_1376F_TAG_SEL_IDX = TAG_SEL_IDX;
											localparam _param_1376F_ARBITER = (CACHE_ENABLE ? "P" : "R");
											localparam _param_1376F_REQ_OUT_BUF = 0;
											localparam _param_1376F_RSP_OUT_BUF = 0;
											if (1) begin : core_bus_nc_arb
												// Trace: src/VX_mem_arb.sv:2:15
												localparam NUM_INPUTS = _param_1376F_NUM_INPUTS;
												// Trace: src/VX_mem_arb.sv:3:15
												localparam NUM_OUTPUTS = _param_1376F_NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:4:15
												localparam DATA_SIZE = _param_1376F_DATA_SIZE;
												// Trace: src/VX_mem_arb.sv:5:15
												localparam TAG_WIDTH = _param_1376F_TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:6:15
												localparam TAG_SEL_IDX = _param_1376F_TAG_SEL_IDX;
												// Trace: src/VX_mem_arb.sv:7:15
												localparam REQ_OUT_BUF = _param_1376F_REQ_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:8:15
												localparam RSP_OUT_BUF = _param_1376F_RSP_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:9:16
												localparam ARBITER = _param_1376F_ARBITER;
												// Trace: src/VX_mem_arb.sv:10:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:11:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_arb.sv:12:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_arb.sv:14:5
												wire clk;
												// Trace: src/VX_mem_arb.sv:15:5
												wire reset;
												// Trace: src/VX_mem_arb.sv:16:5
												localparam _mbase_bus_in_if = 0;
												// Trace: src/VX_mem_arb.sv:17:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_arb.sv:19:5
												localparam DATA_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:20:5
												localparam LOG_NUM_REQS = 0;
												// Trace: src/VX_mem_arb.sv:21:5
												localparam REQ_DATAW = 73;
												// Trace: src/VX_mem_arb.sv:22:5
												localparam RSP_DATAW = 35;
												// Trace: src/VX_mem_arb.sv:24:5
												wire [0:0] req_valid_in;
												// Trace: src/VX_mem_arb.sv:25:5
												wire [72:0] req_data_in;
												// Trace: src/VX_mem_arb.sv:26:5
												wire [0:0] req_ready_in;
												// Trace: src/VX_mem_arb.sv:27:5
												wire [0:0] req_valid_out;
												// Trace: src/VX_mem_arb.sv:28:5
												wire [72:0] req_data_out;
												// Trace: src/VX_mem_arb.sv:29:5
												wire [0:0] req_sel_out;
												// Trace: src/VX_mem_arb.sv:30:5
												wire [0:0] req_ready_out;
												// Trace: src/VX_mem_arb.sv:31:5
												genvar _gv_i_80;
												for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
													localparam i = _gv_i_80;
													// Trace: src/VX_mem_arb.sv:32:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_arb.sv:33:9
													assign req_data_in[i * 73+:73] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_arb.sv:34:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_arb.sv:36:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(REQ_OUT_BUF)
												) req_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(req_valid_in),
													.ready_in(req_ready_in),
													.data_in(req_data_in),
													.data_out(req_data_out),
													.sel_out(req_sel_out),
													.valid_out(req_valid_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_arb.sv:53:5
												genvar _gv_i_81;
												for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
													localparam i = _gv_i_81;
													// Trace: src/VX_mem_arb.sv:54:9
													wire [2:0] req_tag_out;
													// Trace: src/VX_mem_arb.sv:55:9
													VX_bits_insert #(
														.N(TAG_WIDTH),
														.S(LOG_NUM_REQS),
														.POS(TAG_SEL_IDX)
													) bits_insert(
														.data_in(req_tag_out),
														.ins_in(req_sel_out[i+:1]),
														.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[2-:3])
													);
													// Trace: src/VX_mem_arb.sv:64:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_arb.sv:65:9
													assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[72], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[71-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[41-:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[9-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[5-:3], req_tag_out} = req_data_out[i * 73+:73];
													// Trace: src/VX_mem_arb.sv:73:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_ready;
												end
												// Trace: src/VX_mem_arb.sv:75:5
												wire [0:0] rsp_valid_out;
												// Trace: src/VX_mem_arb.sv:76:5
												wire [34:0] rsp_data_out;
												// Trace: src/VX_mem_arb.sv:77:5
												wire [0:0] rsp_ready_out;
												// Trace: src/VX_mem_arb.sv:78:5
												wire [0:0] rsp_valid_in;
												// Trace: src/VX_mem_arb.sv:79:5
												wire [34:0] rsp_data_in;
												// Trace: src/VX_mem_arb.sv:80:5
												wire [0:0] rsp_ready_in;
												// Trace: src/VX_mem_arb.sv:81:5
												if (1) begin : g_passthru
													genvar _gv_i_83;
													for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_83;
														// Trace: src/VX_mem_arb.sv:116:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:117:13
														assign rsp_data_in[i * 35+:35] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_data;
														// Trace: src/VX_mem_arb.sv:118:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:120:9
													VX_stream_arb #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.ARBITER(ARBITER),
														.OUT_BUF(RSP_OUT_BUF)
													) req_arb(
														.clk(clk),
														.reset(reset),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out),
														.sel_out()
													);
												end
												// Trace: src/VX_mem_arb.sv:138:5
												genvar _gv_i_84;
												for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
													localparam i = _gv_i_84;
													// Trace: src/VX_mem_arb.sv:139:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_arb.sv:140:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 35+:35];
													// Trace: src/VX_mem_arb.sv:141:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign core_bus_nc_arb.clk = clk;
											assign core_bus_nc_arb.reset = reset;
											// Trace: src/VX_cache_bypass.sv:102:5
											// expanded interface instance: mem_bus_out_nc_if
											localparam _param_0061C_DATA_SIZE = LINE_SIZE;
											localparam _param_0061C_TAG_WIDTH = MEM_TAG_NC2_WIDTH;
											genvar _arr_0061C;
											for (_arr_0061C = 0; _arr_0061C <= 0; _arr_0061C = _arr_0061C + 1) begin : mem_bus_out_nc_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_0061C_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_0061C_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [612:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [518:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:106:5
											genvar _gv_i_181;
											for (_gv_i_181 = 0; _gv_i_181 < MEM_PORTS; _gv_i_181 = _gv_i_181 + 1) begin : g_mem_bus_out_nc
												localparam i = _gv_i_181;
												// Trace: src/VX_cache_bypass.sv:107:9
												wire core_req_nc_arb_rw;
												// Trace: src/VX_cache_bypass.sv:108:9
												wire [3:0] core_req_nc_arb_byteen;
												// Trace: src/VX_cache_bypass.sv:109:9
												wire [29:0] core_req_nc_arb_addr;
												// Trace: src/VX_cache_bypass.sv:110:9
												wire [2:0] core_req_nc_arb_flags;
												// Trace: src/VX_cache_bypass.sv:111:9
												wire [31:0] core_req_nc_arb_data;
												// Trace: src/VX_cache_bypass.sv:112:9
												wire [2:0] core_req_nc_arb_tag;
												// Trace: src/VX_cache_bypass.sv:113:9
												assign {core_req_nc_arb_rw, core_req_nc_arb_addr, core_req_nc_arb_data, core_req_nc_arb_byteen, core_req_nc_arb_flags, core_req_nc_arb_tag} = core_bus_nc_arb_if[i].req_data;
												// Trace: src/VX_cache_bypass.sv:121:9
												wire [25:0] core_req_nc_arb_addr_w;
												// Trace: src/VX_cache_bypass.sv:122:9
												reg [63:0] core_req_nc_arb_byteen_w;
												// Trace: src/VX_cache_bypass.sv:123:9
												reg [511:0] core_req_nc_arb_data_w;
												// Trace: src/VX_cache_bypass.sv:124:9
												wire [31:0] core_rsp_nc_arb_data_w;
												// Trace: src/VX_cache_bypass.sv:125:9
												wire [6:0] core_req_nc_arb_tag_w;
												// Trace: src/VX_cache_bypass.sv:126:9
												wire [2:0] core_rsp_nc_arb_tag_w;
												if (1) begin : g_multi_word_line
													// Trace: src/VX_cache_bypass.sv:128:13
													wire [3:0] rsp_wsel;
													// Trace: src/VX_cache_bypass.sv:129:13
													wire [3:0] req_wsel = core_req_nc_arb_addr[3:0];
													// Trace: src/VX_cache_bypass.sv:130:13
													always @(*) begin
														// Trace: src/VX_cache_bypass.sv:131:17
														core_req_nc_arb_byteen_w = 1'sb0;
														// Trace: src/VX_cache_bypass.sv:132:17
														core_req_nc_arb_byteen_w[req_wsel * 4+:4] = core_req_nc_arb_byteen;
														// Trace: src/VX_cache_bypass.sv:133:17
														core_req_nc_arb_data_w = 1'sbx;
														// Trace: src/VX_cache_bypass.sv:134:17
														core_req_nc_arb_data_w[req_wsel * 32+:32] = core_req_nc_arb_data;
													end
													// Trace: src/VX_cache_bypass.sv:136:13
													VX_bits_insert #(
														.N(MEM_TAG_NC1_WIDTH),
														.S(WSEL_BITS),
														.POS(TAG_SEL_IDX)
													) wsel_insert(
														.data_in(core_req_nc_arb_tag),
														.ins_in(req_wsel),
														.data_out(core_req_nc_arb_tag_w)
													);
													// Trace: src/VX_cache_bypass.sv:145:13
													VX_bits_remove #(
														.N(MEM_TAG_NC2_WIDTH),
														.S(WSEL_BITS),
														.POS(TAG_SEL_IDX)
													) wsel_remove(
														.data_in(mem_bus_out_nc_if[i].rsp_data[6-:7]),
														.sel_out(rsp_wsel),
														.data_out(core_rsp_nc_arb_tag_w)
													);
													// Trace: src/VX_cache_bypass.sv:154:13
													assign core_req_nc_arb_addr_w = core_req_nc_arb_addr[WSEL_BITS+:MEM_ADDR_WIDTH];
													// Trace: src/VX_cache_bypass.sv:155:13
													assign core_rsp_nc_arb_data_w = mem_bus_out_nc_if[i].rsp_data[7 + (rsp_wsel * CORE_DATA_WIDTH)+:CORE_DATA_WIDTH];
												end
												// Trace: src/VX_cache_bypass.sv:164:9
												assign mem_bus_out_nc_if[i].req_valid = core_bus_nc_arb_if[i].req_valid;
												// Trace: src/VX_cache_bypass.sv:165:9
												assign mem_bus_out_nc_if[i].req_data = {core_req_nc_arb_rw, core_req_nc_arb_addr_w, core_req_nc_arb_data_w, core_req_nc_arb_byteen_w, core_req_nc_arb_flags, core_req_nc_arb_tag_w};
												// Trace: src/VX_cache_bypass.sv:173:9
												assign core_bus_nc_arb_if[i].req_ready = mem_bus_out_nc_if[i].req_ready;
												// Trace: src/VX_cache_bypass.sv:174:9
												assign core_bus_nc_arb_if[i].rsp_valid = mem_bus_out_nc_if[i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:175:9
												assign core_bus_nc_arb_if[i].rsp_data = {core_rsp_nc_arb_data_w, core_rsp_nc_arb_tag_w};
												// Trace: src/VX_cache_bypass.sv:179:9
												assign mem_bus_out_nc_if[i].rsp_ready = core_bus_nc_arb_if[i].rsp_ready;
											end
											// Trace: src/VX_cache_bypass.sv:181:5
											// expanded interface instance: mem_bus_out_src_if
											localparam _param_913F6_DATA_SIZE = LINE_SIZE;
											localparam _param_913F6_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
											genvar _arr_913F6;
											for (_arr_913F6 = 0; _arr_913F6 <= (((CACHE_ENABLE ? 2 : 1) * MEM_PORTS) - 1); _arr_913F6 = _arr_913F6 + 1) begin : mem_bus_out_src_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_913F6_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_913F6_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [612:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [518:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:185:5
											genvar _gv_i_182;
											for (_gv_i_182 = 0; _gv_i_182 < MEM_PORTS; _gv_i_182 = _gv_i_182 + 1) begin : g_mem_bus_out_src
												localparam i = _gv_i_182;
												// Trace: src/VX_cache_bypass.sv:186:5
												assign mem_bus_out_src_if[0 + i].req_valid = mem_bus_out_nc_if[i].req_valid;
												// Trace: src/VX_cache_bypass.sv:187:5
												assign mem_bus_out_src_if[0 + i].req_data[612] = mem_bus_out_nc_if[i].req_data[612];
												// Trace: src/VX_cache_bypass.sv:188:5
												assign mem_bus_out_src_if[0 + i].req_data[611-:26] = mem_bus_out_nc_if[i].req_data[611-:26];
												// Trace: src/VX_cache_bypass.sv:189:5
												assign mem_bus_out_src_if[0 + i].req_data[585-:512] = mem_bus_out_nc_if[i].req_data[585-:512];
												// Trace: src/VX_cache_bypass.sv:190:5
												assign mem_bus_out_src_if[0 + i].req_data[73-:64] = mem_bus_out_nc_if[i].req_data[73-:64];
												// Trace: src/VX_cache_bypass.sv:191:5
												assign mem_bus_out_src_if[0 + i].req_data[9-:3] = mem_bus_out_nc_if[i].req_data[9-:3];
												if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk1
													if (1) begin : genblk1
														if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
															// Trace: src/VX_cache_bypass.sv:196:17
															assign mem_bus_out_src_if[0 + i].req_data[6-:7] = {mem_bus_out_nc_if[i].req_data[6-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_NC2_WIDTH {1'b0}}, mem_bus_out_nc_if[i].req_data[5-:6]};
														end
														else begin : genblk1
															// Trace: src/VX_cache_bypass.sv:198:17
															assign mem_bus_out_src_if[0 + i].req_data[6-:7] = {mem_bus_out_nc_if[i].req_data[6-:1], mem_bus_out_nc_if[i].req_data[(MEM_TAG_OUT_WIDTH - UUID_WIDTH) - 1:0]};
														end
													end
												end
												else begin : genblk1
													// Trace: src/VX_cache_bypass.sv:208:9
													assign mem_bus_out_src_if[0 + i].req_data[6-:7] = mem_bus_out_nc_if[i].req_data[6-:7];
												end
												// Trace: src/VX_cache_bypass.sv:211:5
												assign mem_bus_out_nc_if[i].req_ready = mem_bus_out_src_if[0 + i].req_ready;
												// Trace: src/VX_cache_bypass.sv:212:5
												assign mem_bus_out_nc_if[i].rsp_valid = mem_bus_out_src_if[0 + i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:213:5
												assign mem_bus_out_nc_if[i].rsp_data[518-:512] = mem_bus_out_src_if[0 + i].rsp_data[518-:512];
												if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk2
													if (1) begin : genblk1
														if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
															// Trace: src/VX_cache_bypass.sv:218:17
															assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[6-:1], mem_bus_out_src_if[0 + i].rsp_data[5:0]};
														end
														else begin : genblk1
															// Trace: src/VX_cache_bypass.sv:220:17
															assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[6-:1], {MEM_TAG_NC2_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[0 + i].rsp_data[5-:6]};
														end
													end
												end
												else begin : genblk2
													// Trace: src/VX_cache_bypass.sv:230:9
													assign mem_bus_out_nc_if[i].rsp_data[6-:7] = mem_bus_out_src_if[0 + i].rsp_data[6-:7];
												end
												// Trace: src/VX_cache_bypass.sv:233:5
												assign mem_bus_out_src_if[0 + i].rsp_ready = mem_bus_out_nc_if[i].rsp_ready;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:235:5
													assign mem_bus_out_src_if[1 + i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_valid;
													// Trace: src/VX_cache_bypass.sv:236:5
													assign mem_bus_out_src_if[1 + i].req_data[612] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[610];
													// Trace: src/VX_cache_bypass.sv:237:5
													assign mem_bus_out_src_if[1 + i].req_data[611-:26] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[609-:26];
													// Trace: src/VX_cache_bypass.sv:238:5
													assign mem_bus_out_src_if[1 + i].req_data[585-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[583-:512];
													// Trace: src/VX_cache_bypass.sv:239:5
													assign mem_bus_out_src_if[1 + i].req_data[73-:64] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[71-:64];
													// Trace: src/VX_cache_bypass.sv:240:5
													assign mem_bus_out_src_if[1 + i].req_data[9-:3] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[7-:3];
													if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk1
														if (1) begin : genblk1
															if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
																// Trace: src/VX_cache_bypass.sv:245:17
																assign mem_bus_out_src_if[1 + i].req_data[6-:7] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_IN_WIDTH {1'b0}}, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[3-:4]};
															end
															else begin : genblk1
																// Trace: src/VX_cache_bypass.sv:247:17
																assign mem_bus_out_src_if[1 + i].req_data[6-:7] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[(MEM_TAG_OUT_WIDTH - UUID_WIDTH) - 1:0]};
															end
														end
													end
													else begin : genblk1
														// Trace: src/VX_cache_bypass.sv:257:9
														assign mem_bus_out_src_if[1 + i].req_data[6-:7] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:5];
													end
													// Trace: src/VX_cache_bypass.sv:260:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = mem_bus_out_src_if[1 + i].req_ready;
													// Trace: src/VX_cache_bypass.sv:261:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = mem_bus_out_src_if[1 + i].rsp_valid;
													// Trace: src/VX_cache_bypass.sv:262:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[516-:512] = mem_bus_out_src_if[1 + i].rsp_data[518-:512];
													if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk2
														if (1) begin : genblk1
															if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
																// Trace: src/VX_cache_bypass.sv:267:17
																assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[6-:1], mem_bus_out_src_if[1 + i].rsp_data[3:0]};
															end
															else begin : genblk1
																// Trace: src/VX_cache_bypass.sv:269:17
																assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[6-:1], {MEM_TAG_IN_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[1 + i].rsp_data[5-:6]};
															end
														end
													end
													else begin : genblk2
														// Trace: src/VX_cache_bypass.sv:279:9
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = mem_bus_out_src_if[1 + i].rsp_data[6-:7];
													end
													// Trace: src/VX_cache_bypass.sv:282:5
													assign mem_bus_out_src_if[1 + i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_ready;
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:284:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = 0;
													// Trace: src/VX_cache_bypass.sv:285:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = 0;
													// Trace: src/VX_cache_bypass.sv:286:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data = 1'sb0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:289:5
											// expanded module instance: mem_bus_out_arb
											localparam _bbase_B06D0_bus_in_if = 0;
											localparam _bbase_B06D0_bus_out_if = 0;
											localparam _param_B06D0_NUM_INPUTS = (CACHE_ENABLE ? 2 : 1) * MEM_PORTS;
											localparam _param_B06D0_NUM_OUTPUTS = MEM_PORTS;
											localparam _param_B06D0_DATA_SIZE = LINE_SIZE;
											localparam _param_B06D0_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
											localparam _param_B06D0_ARBITER = "R";
											localparam _param_B06D0_REQ_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
											localparam _param_B06D0_RSP_OUT_BUF = 0;
											if (1) begin : mem_bus_out_arb
												// Trace: src/VX_mem_arb.sv:2:15
												localparam NUM_INPUTS = _param_B06D0_NUM_INPUTS;
												// Trace: src/VX_mem_arb.sv:3:15
												localparam NUM_OUTPUTS = _param_B06D0_NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:4:15
												localparam DATA_SIZE = _param_B06D0_DATA_SIZE;
												// Trace: src/VX_mem_arb.sv:5:15
												localparam TAG_WIDTH = _param_B06D0_TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:6:15
												localparam TAG_SEL_IDX = 0;
												// Trace: src/VX_mem_arb.sv:7:15
												localparam REQ_OUT_BUF = _param_B06D0_REQ_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:8:15
												localparam RSP_OUT_BUF = _param_B06D0_RSP_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:9:16
												localparam ARBITER = _param_B06D0_ARBITER;
												// Trace: src/VX_mem_arb.sv:10:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:11:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_arb.sv:12:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_arb.sv:14:5
												wire clk;
												// Trace: src/VX_mem_arb.sv:15:5
												wire reset;
												// Trace: src/VX_mem_arb.sv:16:5
												localparam _mbase_bus_in_if = 0;
												// Trace: src/VX_mem_arb.sv:17:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_arb.sv:19:5
												localparam DATA_WIDTH = 512;
												// Trace: src/VX_mem_arb.sv:20:5
												localparam LOG_NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? $clog2((NUM_INPUTS + 0) / 1) : 0);
												// Trace: src/VX_mem_arb.sv:21:5
												localparam REQ_DATAW = 606 + TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:22:5
												localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:24:5
												wire [NUM_INPUTS - 1:0] req_valid_in;
												// Trace: src/VX_mem_arb.sv:25:5
												wire [(NUM_INPUTS * REQ_DATAW) - 1:0] req_data_in;
												// Trace: src/VX_mem_arb.sv:26:5
												wire [NUM_INPUTS - 1:0] req_ready_in;
												// Trace: src/VX_mem_arb.sv:27:5
												wire [0:0] req_valid_out;
												// Trace: src/VX_mem_arb.sv:28:5
												wire [REQ_DATAW - 1:0] req_data_out;
												// Trace: src/VX_mem_arb.sv:29:5
												wire [(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1) - 1:0] req_sel_out;
												// Trace: src/VX_mem_arb.sv:30:5
												wire [0:0] req_ready_out;
												// Trace: src/VX_mem_arb.sv:31:5
												genvar _gv_i_80;
												for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
													localparam i = _gv_i_80;
													// Trace: src/VX_mem_arb.sv:32:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_arb.sv:33:9
													assign req_data_in[i * 613+:613] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_arb.sv:34:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_arb.sv:36:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(REQ_OUT_BUF)
												) req_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(req_valid_in),
													.ready_in(req_ready_in),
													.data_in(req_data_in),
													.data_out(req_data_out),
													.sel_out(req_sel_out),
													.valid_out(req_valid_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_arb.sv:53:5
												genvar _gv_i_81;
												for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
													localparam i = _gv_i_81;
													// Trace: src/VX_mem_arb.sv:54:9
													wire [TAG_WIDTH - 1:0] req_tag_out;
													// Trace: src/VX_mem_arb.sv:55:9
													VX_bits_insert #(
														.N(TAG_WIDTH),
														.S(LOG_NUM_REQS),
														.POS(TAG_SEL_IDX)
													) bits_insert(
														.data_in(req_tag_out),
														.ins_in(req_sel_out[i * 1+:1]),
														.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[4-:5])
													);
													// Trace: src/VX_mem_arb.sv:64:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_arb.sv:65:9
													assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[610], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[609-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[583-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[71-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[7-:3], req_tag_out} = req_data_out[i * 613+:613];
													// Trace: src/VX_mem_arb.sv:73:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
												end
												// Trace: src/VX_mem_arb.sv:75:5
												wire [NUM_INPUTS - 1:0] rsp_valid_out;
												// Trace: src/VX_mem_arb.sv:76:5
												wire [(NUM_INPUTS * RSP_DATAW) - 1:0] rsp_data_out;
												// Trace: src/VX_mem_arb.sv:77:5
												wire [NUM_INPUTS - 1:0] rsp_ready_out;
												// Trace: src/VX_mem_arb.sv:78:5
												wire [0:0] rsp_valid_in;
												// Trace: src/VX_mem_arb.sv:79:5
												wire [RSP_DATAW - 1:0] rsp_data_in;
												// Trace: src/VX_mem_arb.sv:80:5
												wire [0:0] rsp_ready_in;
												// Trace: src/VX_mem_arb.sv:81:5
												if (NUM_INPUTS > NUM_OUTPUTS) begin : g_rsp_enabled
													// Trace: src/VX_mem_arb.sv:82:9
													wire [LOG_NUM_REQS - 1:0] rsp_sel_in;
													genvar _gv_i_82;
													for (_gv_i_82 = 0; _gv_i_82 < NUM_OUTPUTS; _gv_i_82 = _gv_i_82 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_82;
														// Trace: src/VX_mem_arb.sv:84:13
														wire [TAG_WIDTH - 1:0] rsp_tag_out;
														// Trace: src/VX_mem_arb.sv:85:13
														VX_bits_remove #(
															.N(TAG_WIDTH + LOG_NUM_REQS),
															.S(LOG_NUM_REQS),
															.POS(TAG_SEL_IDX)
														) bits_remove(
															.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[4-:5]),
															.sel_out(rsp_sel_in[i * 1+:1]),
															.data_out(rsp_tag_out)
														);
														// Trace: src/VX_mem_arb.sv:94:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:95:13
														assign rsp_data_in[i * 519+:519] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[516-:512], rsp_tag_out};
														// Trace: src/VX_mem_arb.sv:96:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:98:9
													VX_stream_switch #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.OUT_BUF(RSP_OUT_BUF)
													) rsp_switch(
														.clk(clk),
														.reset(reset),
														.sel_in(rsp_sel_in),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out)
													);
												end
												else begin : g_passthru
													genvar _gv_i_83;
													for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_83;
														// Trace: src/VX_mem_arb.sv:116:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:117:13
														assign rsp_data_in[i * 519+:519] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
														// Trace: src/VX_mem_arb.sv:118:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:120:9
													VX_stream_arb #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.ARBITER(ARBITER),
														.OUT_BUF(RSP_OUT_BUF)
													) req_arb(
														.clk(clk),
														.reset(reset),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out),
														.sel_out()
													);
												end
												// Trace: src/VX_mem_arb.sv:138:5
												genvar _gv_i_84;
												for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
													localparam i = _gv_i_84;
													// Trace: src/VX_mem_arb.sv:139:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_arb.sv:140:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
													// Trace: src/VX_mem_arb.sv:141:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign mem_bus_out_arb.clk = clk;
											assign mem_bus_out_arb.reset = reset;
										end
										assign cache_bypass.clk = clk;
										assign cache_bypass.reset = reset;
									end
									else begin : g_no_bypass
										genvar _gv_i_167;
										for (_gv_i_167 = 0; _gv_i_167 < NUM_REQS; _gv_i_167 = _gv_i_167 + 1) begin : g_core_bus_cache_if
											localparam i = _gv_i_167;
											// Trace: src/VX_cache_wrap.sv:76:5
											assign core_bus_cache_if[i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].req_valid;
											// Trace: src/VX_cache_wrap.sv:77:5
											assign core_bus_cache_if[i].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].req_data;
											// Trace: src/VX_cache_wrap.sv:78:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].req_ready = core_bus_cache_if[i].req_ready;
											// Trace: src/VX_cache_wrap.sv:79:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_valid = core_bus_cache_if[i].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:80:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_data = core_bus_cache_if[i].rsp_data;
											// Trace: src/VX_cache_wrap.sv:81:5
											assign core_bus_cache_if[i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_ready;
										end
										genvar _gv_i_168;
										for (_gv_i_168 = 0; _gv_i_168 < MEM_PORTS; _gv_i_168 = _gv_i_168 + 1) begin : g_mem_bus_tmp_if
											localparam i = _gv_i_168;
											// Trace: src/VX_cache_wrap.sv:84:5
											assign mem_bus_tmp_if[i].req_valid = mem_bus_cache_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:85:5
											assign mem_bus_tmp_if[i].req_data = mem_bus_cache_if[i].req_data;
											// Trace: src/VX_cache_wrap.sv:86:5
											assign mem_bus_cache_if[i].req_ready = mem_bus_tmp_if[i].req_ready;
											// Trace: src/VX_cache_wrap.sv:87:5
											assign mem_bus_cache_if[i].rsp_valid = mem_bus_tmp_if[i].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:88:5
											assign mem_bus_cache_if[i].rsp_data = mem_bus_tmp_if[i].rsp_data;
											// Trace: src/VX_cache_wrap.sv:89:5
											assign mem_bus_tmp_if[i].rsp_ready = mem_bus_cache_if[i].rsp_ready;
										end
									end
									// Trace: src/VX_cache_wrap.sv:92:5
									genvar _gv_i_169;
									for (_gv_i_169 = 0; _gv_i_169 < MEM_PORTS; _gv_i_169 = _gv_i_169 + 1) begin : g_mem_bus_if
										localparam i = _gv_i_169;
										if (WRITE_ENABLE) begin : g_we
											// Trace: src/VX_cache_wrap.sv:94:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:95:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
											// Trace: src/VX_cache_wrap.sv:96:5
											assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
											// Trace: src/VX_cache_wrap.sv:97:5
											assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:98:5
											assign mem_bus_tmp_if[i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
											// Trace: src/VX_cache_wrap.sv:99:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
										end
										else begin : g_ro
											// Trace: src/VX_cache_wrap.sv:101:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:102:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[610] = 0;
											// Trace: src/VX_cache_wrap.sv:103:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[609-:26] = mem_bus_tmp_if[i].req_data[609-:26];
											// Trace: src/VX_cache_wrap.sv:104:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[583-:512] = 1'sb0;
											// Trace: src/VX_cache_wrap.sv:105:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[71-:64] = 1'sb1;
											// Trace: src/VX_cache_wrap.sv:106:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[7-:3] = mem_bus_tmp_if[i].req_data[7-:3];
											// Trace: src/VX_cache_wrap.sv:107:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[4-:5] = mem_bus_tmp_if[i].req_data[4-:5];
											// Trace: src/VX_cache_wrap.sv:108:5
											assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
											// Trace: src/VX_cache_wrap.sv:109:5
											assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:110:5
											assign mem_bus_tmp_if[i].rsp_data[516-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[516-:512];
											// Trace: src/VX_cache_wrap.sv:111:5
											assign mem_bus_tmp_if[i].rsp_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[4-:5];
											// Trace: src/VX_cache_wrap.sv:112:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
										end
									end
									// Trace: src/VX_cache_wrap.sv:115:5
									if (1) begin : g_cache
										// Trace: src/VX_cache_wrap.sv:116:9
										// expanded module instance: cache
										localparam _bbase_90EE2_core_bus_if = 0;
										localparam _bbase_90EE2_mem_bus_if = 0;
										localparam _param_90EE2_INSTANCE_ID = INSTANCE_ID;
										localparam _param_90EE2_CACHE_SIZE = CACHE_SIZE;
										localparam _param_90EE2_LINE_SIZE = LINE_SIZE;
										localparam _param_90EE2_NUM_BANKS = NUM_BANKS;
										localparam _param_90EE2_NUM_WAYS = NUM_WAYS;
										localparam _param_90EE2_WORD_SIZE = WORD_SIZE;
										localparam _param_90EE2_NUM_REQS = NUM_REQS;
										localparam _param_90EE2_MEM_PORTS = MEM_PORTS;
										localparam _param_90EE2_WRITE_ENABLE = WRITE_ENABLE;
										localparam _param_90EE2_WRITEBACK = WRITEBACK;
										localparam _param_90EE2_DIRTY_BYTES = DIRTY_BYTES;
										localparam _param_90EE2_REPL_POLICY = REPL_POLICY;
										localparam _param_90EE2_CRSQ_SIZE = CRSQ_SIZE;
										localparam _param_90EE2_MSHR_SIZE = MSHR_SIZE;
										localparam _param_90EE2_MRSQ_SIZE = MRSQ_SIZE;
										localparam _param_90EE2_MREQ_SIZE = MREQ_SIZE;
										localparam _param_90EE2_UUID_WIDTH = UUID_WIDTH;
										localparam _param_90EE2_TAG_WIDTH = TAG_WIDTH;
										localparam _param_90EE2_FLAGS_WIDTH = FLAGS_WIDTH;
										localparam _param_90EE2_CORE_OUT_BUF = (BYPASS_ENABLE ? 1 : CORE_OUT_BUF);
										localparam _param_90EE2_MEM_OUT_BUF = (BYPASS_ENABLE ? 1 : MEM_OUT_BUF);
										if (1) begin : cache
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_cache.sv:2:16
											localparam INSTANCE_ID = _param_90EE2_INSTANCE_ID;
											// Trace: src/VX_cache.sv:3:15
											localparam NUM_REQS = _param_90EE2_NUM_REQS;
											// Trace: src/VX_cache.sv:4:15
											localparam MEM_PORTS = _param_90EE2_MEM_PORTS;
											// Trace: src/VX_cache.sv:5:15
											localparam CACHE_SIZE = _param_90EE2_CACHE_SIZE;
											// Trace: src/VX_cache.sv:6:15
											localparam LINE_SIZE = _param_90EE2_LINE_SIZE;
											// Trace: src/VX_cache.sv:7:15
											localparam NUM_BANKS = _param_90EE2_NUM_BANKS;
											// Trace: src/VX_cache.sv:8:15
											localparam NUM_WAYS = _param_90EE2_NUM_WAYS;
											// Trace: src/VX_cache.sv:9:15
											localparam WORD_SIZE = _param_90EE2_WORD_SIZE;
											// Trace: src/VX_cache.sv:10:15
											localparam CRSQ_SIZE = _param_90EE2_CRSQ_SIZE;
											// Trace: src/VX_cache.sv:11:15
											localparam MSHR_SIZE = _param_90EE2_MSHR_SIZE;
											// Trace: src/VX_cache.sv:12:15
											localparam MRSQ_SIZE = _param_90EE2_MRSQ_SIZE;
											// Trace: src/VX_cache.sv:13:15
											localparam MREQ_SIZE = _param_90EE2_MREQ_SIZE;
											// Trace: src/VX_cache.sv:14:15
											localparam WRITE_ENABLE = _param_90EE2_WRITE_ENABLE;
											// Trace: src/VX_cache.sv:15:15
											localparam WRITEBACK = _param_90EE2_WRITEBACK;
											// Trace: src/VX_cache.sv:16:15
											localparam DIRTY_BYTES = _param_90EE2_DIRTY_BYTES;
											// Trace: src/VX_cache.sv:17:15
											localparam REPL_POLICY = _param_90EE2_REPL_POLICY;
											// Trace: src/VX_cache.sv:18:15
											localparam UUID_WIDTH = _param_90EE2_UUID_WIDTH;
											// Trace: src/VX_cache.sv:19:15
											localparam TAG_WIDTH = _param_90EE2_TAG_WIDTH;
											// Trace: src/VX_cache.sv:20:15
											localparam FLAGS_WIDTH = _param_90EE2_FLAGS_WIDTH;
											// Trace: src/VX_cache.sv:21:15
											localparam CORE_OUT_BUF = _param_90EE2_CORE_OUT_BUF;
											// Trace: src/VX_cache.sv:22:15
											localparam MEM_OUT_BUF = _param_90EE2_MEM_OUT_BUF;
											// Trace: src/VX_cache.sv:24:5
											wire clk;
											// Trace: src/VX_cache.sv:25:5
											wire reset;
											// Trace: src/VX_cache.sv:26:5
											localparam _mbase_core_bus_if = 0;
											// Trace: src/VX_cache.sv:27:5
											localparam _mbase_mem_bus_if = 0;
											// Trace: src/VX_cache.sv:29:5
											localparam REQ_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:30:5
											localparam WORD_SEL_WIDTH = 4;
											// Trace: src/VX_cache.sv:31:5
											localparam MSHR_ADDR_WIDTH = 4;
											// Trace: src/VX_cache.sv:32:5
											localparam MEM_TAG_WIDTH = 5;
											// Trace: src/VX_cache.sv:34:5
											localparam WORDS_PER_LINE = 16;
											// Trace: src/VX_cache.sv:35:5
											localparam WORD_WIDTH = 32;
											// Trace: src/VX_cache.sv:36:5
											localparam WORD_SEL_BITS = 4;
											// Trace: src/VX_cache.sv:37:5
											localparam BANK_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:38:5
											localparam BANK_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:39:5
											localparam LINE_ADDR_WIDTH = 26;
											// Trace: src/VX_cache.sv:40:5
											localparam CORE_REQ_DATAW = 71;
											// Trace: src/VX_cache.sv:41:5
											localparam CORE_RSP_DATAW = 35;
											// Trace: src/VX_cache.sv:42:5
											localparam BANK_MEM_TAG_WIDTH = 5;
											// Trace: src/VX_cache.sv:43:5
											localparam MEM_REQ_DATAW = 609;
											// Trace: src/VX_cache.sv:44:5
											localparam MEM_RSP_DATAW = 517;
											// Trace: src/VX_cache.sv:45:5
											localparam MEM_PORTS_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:46:5
											localparam MEM_PORTS_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:47:5
											localparam MEM_ARB_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:48:5
											localparam MEM_ARB_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:49:5
											localparam CORE_RSP_REG_DISABLE = 1'd0;
											// Trace: src/VX_cache.sv:50:5
											localparam MEM_REQ_REG_DISABLE = 1'd0;
											// Trace: src/VX_cache.sv:51:5
											localparam REQ_XBAR_BUF = 0;
											// Trace: src/VX_cache.sv:52:5
											// expanded interface instance: core_bus2_if
											localparam _param_9260A_DATA_SIZE = WORD_SIZE;
											localparam _param_9260A_TAG_WIDTH = TAG_WIDTH;
											genvar _arr_9260A;
											for (_arr_9260A = 0; _arr_9260A <= 0; _arr_9260A = _arr_9260A + 1) begin : core_bus2_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_9260A_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_9260A_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [72:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [34:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache.sv:56:5
											wire [0:0] per_bank_flush_begin;
											// Trace: src/VX_cache.sv:57:5
											wire [0:0] flush_uuid;
											// Trace: src/VX_cache.sv:58:5
											wire [0:0] per_bank_flush_end;
											// Trace: src/VX_cache.sv:59:5
											wire [0:0] per_bank_core_req_fire;
											// Trace: src/VX_cache.sv:60:5
											// expanded module instance: flush_unit
											localparam _bbase_1DACF_core_bus_in_if = 0;
											localparam _bbase_1DACF_core_bus_out_if = 0;
											localparam _param_1DACF_NUM_REQS = NUM_REQS;
											localparam _param_1DACF_NUM_BANKS = NUM_BANKS;
											localparam _param_1DACF_UUID_WIDTH = UUID_WIDTH;
											localparam _param_1DACF_TAG_WIDTH = TAG_WIDTH;
											localparam _param_1DACF_BANK_SEL_LATENCY = 0;
											if (1) begin : flush_unit
												// Trace: src/VX_cache_flush.sv:2:15
												localparam NUM_REQS = _param_1DACF_NUM_REQS;
												// Trace: src/VX_cache_flush.sv:3:15
												localparam NUM_BANKS = _param_1DACF_NUM_BANKS;
												// Trace: src/VX_cache_flush.sv:4:15
												localparam UUID_WIDTH = _param_1DACF_UUID_WIDTH;
												// Trace: src/VX_cache_flush.sv:5:15
												localparam TAG_WIDTH = _param_1DACF_TAG_WIDTH;
												// Trace: src/VX_cache_flush.sv:6:15
												localparam BANK_SEL_LATENCY = _param_1DACF_BANK_SEL_LATENCY;
												// Trace: src/VX_cache_flush.sv:8:5
												wire clk;
												// Trace: src/VX_cache_flush.sv:9:5
												wire reset;
												// Trace: src/VX_cache_flush.sv:10:5
												localparam _mbase_core_bus_in_if = 0;
												// Trace: src/VX_cache_flush.sv:11:5
												localparam _mbase_core_bus_out_if = 0;
												// Trace: src/VX_cache_flush.sv:12:5
												wire [0:0] bank_req_fire;
												// Trace: src/VX_cache_flush.sv:13:5
												wire [0:0] flush_begin;
												// Trace: src/VX_cache_flush.sv:14:5
												wire [0:0] flush_uuid;
												// Trace: src/VX_cache_flush.sv:15:5
												wire [0:0] flush_end;
												// Trace: src/VX_cache_flush.sv:17:5
												localparam STATE_IDLE = 0;
												// Trace: src/VX_cache_flush.sv:18:5
												localparam STATE_WAIT1 = 1;
												// Trace: src/VX_cache_flush.sv:19:5
												localparam STATE_FLUSH = 2;
												// Trace: src/VX_cache_flush.sv:20:5
												localparam STATE_WAIT2 = 3;
												// Trace: src/VX_cache_flush.sv:21:5
												localparam STATE_DONE = 4;
												// Trace: src/VX_cache_flush.sv:22:5
												reg [2:0] state;
												reg [2:0] state_n;
												// Trace: src/VX_cache_flush.sv:23:5
												wire no_inflight_reqs;
												// Trace: src/VX_cache_flush.sv:24:5
												if (1) begin : g_no_bank_sel_latency
													// Trace: src/VX_cache_flush.sv:63:9
													assign no_inflight_reqs = 0;
												end
												// Trace: src/VX_cache_flush.sv:65:5
												reg [0:0] flush_done;
												reg [0:0] flush_done_n;
												// Trace: src/VX_cache_flush.sv:66:5
												wire [0:0] flush_req_mask;
												// Trace: src/VX_cache_flush.sv:67:5
												genvar _gv_i_116;
												for (_gv_i_116 = 0; _gv_i_116 < NUM_REQS; _gv_i_116 = _gv_i_116 + 1) begin : g_flush_req_mask
													localparam i = _gv_i_116;
													// Trace: src/VX_cache_flush.sv:68:9
													assign flush_req_mask[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data[3];
												end
												// Trace: src/VX_cache_flush.sv:70:5
												wire flush_req_enable = |flush_req_mask;
												// Trace: src/VX_cache_flush.sv:71:5
												reg [0:0] lock_released;
												reg [0:0] lock_released_n;
												// Trace: src/VX_cache_flush.sv:72:5
												reg [0:0] flush_uuid_r;
												reg [0:0] flush_uuid_n;
												// Trace: src/VX_cache_flush.sv:73:5
												genvar _gv_i_117;
												for (_gv_i_117 = 0; _gv_i_117 < NUM_REQS; _gv_i_117 = _gv_i_117 + 1) begin : g_core_bus_out_req
													localparam i = _gv_i_117;
													// Trace: src/VX_cache_flush.sv:74:9
													wire input_enable = ~flush_req_enable || lock_released[i];
													// Trace: src/VX_cache_flush.sv:75:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_valid && input_enable;
													// Trace: src/VX_cache_flush.sv:76:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data;
													// Trace: src/VX_cache_flush.sv:77:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_ready && input_enable;
												end
												// Trace: src/VX_cache_flush.sv:79:5
												genvar _gv_i_118;
												for (_gv_i_118 = 0; _gv_i_118 < NUM_REQS; _gv_i_118 = _gv_i_118 + 1) begin : g_core_bus_in_rsp
													localparam i = _gv_i_118;
													// Trace: src/VX_cache_flush.sv:80:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_valid;
													// Trace: src/VX_cache_flush.sv:81:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_data;
													// Trace: src/VX_cache_flush.sv:82:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_ready;
												end
												// Trace: src/VX_cache_flush.sv:84:5
												reg [0:0] core_bus_out_uuid;
												// Trace: src/VX_cache_flush.sv:85:5
												wire [0:0] core_bus_out_ready;
												// Trace: src/VX_cache_flush.sv:86:5
												genvar _gv_i_119;
												for (_gv_i_119 = 0; _gv_i_119 < NUM_REQS; _gv_i_119 = _gv_i_119 + 1) begin : g_core_bus_out_uuid
													localparam i = _gv_i_119;
													if (1) begin : g_uuid
														// Trace: src/VX_cache_flush.sv:88:13
														wire [1:1] sv2v_tmp_F411A;
														assign sv2v_tmp_F411A = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data[2-:1];
														always @(*) core_bus_out_uuid[i+:1] = sv2v_tmp_F411A;
													end
												end
												// Trace: src/VX_cache_flush.sv:93:5
												genvar _gv_i_120;
												for (_gv_i_120 = 0; _gv_i_120 < NUM_REQS; _gv_i_120 = _gv_i_120 + 1) begin : g_core_bus_out_ready
													localparam i = _gv_i_120;
													// Trace: src/VX_cache_flush.sv:94:9
													assign core_bus_out_ready[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_ready;
												end
												// Trace: src/VX_cache_flush.sv:96:5
												always @(*) begin
													// Trace: src/VX_cache_flush.sv:97:9
													state_n = state;
													// Trace: src/VX_cache_flush.sv:98:9
													flush_done_n = flush_done;
													// Trace: src/VX_cache_flush.sv:99:9
													lock_released_n = lock_released;
													// Trace: src/VX_cache_flush.sv:100:9
													flush_uuid_n = flush_uuid_r;
													// Trace: src/VX_cache_flush.sv:101:9
													case (state)
														default:
															// Trace: src/VX_cache_flush.sv:103:17
															if (flush_req_enable) begin
																// Trace: src/VX_cache_flush.sv:104:21
																state_n = STATE_FLUSH;
																// Trace: src/VX_cache_flush.sv:105:21
																begin : sv2v_autoblock_1
																	// Trace: src/VX_cache_flush.sv:105:26
																	integer i;
																	// Trace: src/VX_cache_flush.sv:105:26
																	for (i = 0; i >= 0; i = i - 1)
																		begin
																			// Trace: src/VX_cache_flush.sv:106:25
																			if (flush_req_mask[i])
																				// Trace: src/VX_cache_flush.sv:107:29
																				flush_uuid_n = core_bus_out_uuid[i+:1];
																		end
																end
															end
														STATE_WAIT1:
															// Trace: src/VX_cache_flush.sv:113:17
															if (no_inflight_reqs)
																// Trace: src/VX_cache_flush.sv:114:21
																state_n = STATE_FLUSH;
														STATE_FLUSH:
															// Trace: src/VX_cache_flush.sv:118:17
															state_n = STATE_WAIT2;
														STATE_WAIT2: begin
															// Trace: src/VX_cache_flush.sv:121:17
															flush_done_n = flush_done | flush_end;
															// Trace: src/VX_cache_flush.sv:122:17
															if (flush_done_n == {NUM_BANKS {1'b1}}) begin
																// Trace: src/VX_cache_flush.sv:123:21
																state_n = STATE_DONE;
																// Trace: src/VX_cache_flush.sv:124:21
																flush_done_n = 1'sb0;
																// Trace: src/VX_cache_flush.sv:125:21
																lock_released_n = flush_req_mask;
															end
														end
														STATE_DONE: begin
															// Trace: src/VX_cache_flush.sv:129:17
															lock_released_n = lock_released & ~core_bus_out_ready;
															// Trace: src/VX_cache_flush.sv:130:17
															if (lock_released_n == 0)
																// Trace: src/VX_cache_flush.sv:131:21
																state_n = STATE_IDLE;
														end
													endcase
												end
												// Trace: src/VX_cache_flush.sv:136:5
												always @(posedge clk) begin
													// Trace: src/VX_cache_flush.sv:137:9
													if (reset) begin
														// Trace: src/VX_cache_flush.sv:138:13
														state <= STATE_IDLE;
														// Trace: src/VX_cache_flush.sv:139:13
														flush_done <= 1'sb0;
														// Trace: src/VX_cache_flush.sv:140:13
														lock_released <= 1'sb0;
													end
													else begin
														// Trace: src/VX_cache_flush.sv:142:13
														state <= state_n;
														// Trace: src/VX_cache_flush.sv:143:13
														flush_done <= flush_done_n;
														// Trace: src/VX_cache_flush.sv:144:13
														lock_released <= lock_released_n;
													end
													// Trace: src/VX_cache_flush.sv:146:9
													flush_uuid_r <= flush_uuid_n;
												end
												// Trace: src/VX_cache_flush.sv:148:5
												assign flush_begin = {NUM_BANKS {state == STATE_FLUSH}};
												// Trace: src/VX_cache_flush.sv:149:5
												assign flush_uuid = flush_uuid_r;
											end
											assign flush_unit.clk = clk;
											assign flush_unit.reset = reset;
											assign flush_unit.bank_req_fire = per_bank_core_req_fire;
											assign per_bank_flush_begin = flush_unit.flush_begin;
											assign flush_uuid = flush_unit.flush_uuid;
											assign flush_unit.flush_end = per_bank_flush_end;
											// Trace: src/VX_cache.sv:76:5
											// expanded interface instance: mem_bus_tmp_if
											localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
											localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
											genvar _arr_4FE36;
											for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [610:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [516:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache.sv:80:5
											wire [0:0] mem_rsp_queue_valid;
											// Trace: src/VX_cache.sv:81:5
											wire [516:0] mem_rsp_queue_data;
											// Trace: src/VX_cache.sv:82:5
											wire [0:0] mem_rsp_queue_ready;
											// Trace: src/VX_cache.sv:83:5
											genvar _gv_i_29;
											for (_gv_i_29 = 0; _gv_i_29 < MEM_PORTS; _gv_i_29 = _gv_i_29 + 1) begin : g_mem_rsp_queue
												localparam i = _gv_i_29;
												// Trace: src/VX_cache.sv:84:9
												VX_elastic_buffer #(
													.DATAW(MEM_RSP_DATAW),
													.SIZE(MRSQ_SIZE),
													.OUT_REG(1'd0)
												) mem_rsp_queue(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_bus_tmp_if[i].rsp_valid),
													.data_in(mem_bus_tmp_if[i].rsp_data),
													.ready_in(mem_bus_tmp_if[i].rsp_ready),
													.valid_out(mem_rsp_queue_valid[i]),
													.data_out(mem_rsp_queue_data[i * 517+:517]),
													.ready_out(mem_rsp_queue_ready[i])
												);
											end
											// Trace: src/VX_cache.sv:99:5
											wire [516:0] mem_rsp_queue_data_s;
											// Trace: src/VX_cache.sv:100:5
											wire [0:0] mem_rsp_queue_sel;
											// Trace: src/VX_cache.sv:101:5
											genvar _gv_i_30;
											for (_gv_i_30 = 0; _gv_i_30 < MEM_PORTS; _gv_i_30 = _gv_i_30 + 1) begin : g_mem_rsp_queue_data_s
												localparam i = _gv_i_30;
												// Trace: src/VX_cache.sv:102:9
												wire [4:0] mem_rsp_tag_s = mem_rsp_queue_data[(i * 517) + 4-:5];
												// Trace: src/VX_cache.sv:103:9
												wire [511:0] mem_rsp_data_s = mem_rsp_queue_data[(i * 517) + 516-:512];
												// Trace: src/VX_cache.sv:104:9
												assign mem_rsp_queue_data_s[i * 517+:517] = {mem_rsp_data_s, mem_rsp_tag_s};
											end
											// Trace: src/VX_cache.sv:106:5
											genvar _gv_i_31;
											for (_gv_i_31 = 0; _gv_i_31 < MEM_PORTS; _gv_i_31 = _gv_i_31 + 1) begin : g_mem_rsp_queue_sel
												localparam i = _gv_i_31;
												if (1) begin : g_singlebank
													// Trace: src/VX_cache.sv:121:13
													assign mem_rsp_queue_sel[i+:1] = 0;
												end
											end
											// Trace: src/VX_cache.sv:124:5
											wire [0:0] per_bank_mem_rsp_valid;
											// Trace: src/VX_cache.sv:125:5
											wire [516:0] per_bank_mem_rsp_pdata;
											// Trace: src/VX_cache.sv:126:5
											wire [0:0] per_bank_mem_rsp_ready;
											// Trace: src/VX_cache.sv:127:5
											VX_stream_omega #(
												.NUM_INPUTS(MEM_PORTS),
												.NUM_OUTPUTS(NUM_BANKS),
												.DATAW(517),
												.ARBITER("R"),
												.OUT_BUF(3)
											) mem_rsp_xbar(
												.clk(clk),
												.reset(reset),
												.valid_in(mem_rsp_queue_valid),
												.data_in(mem_rsp_queue_data_s),
												.sel_in(mem_rsp_queue_sel),
												.ready_in(mem_rsp_queue_ready),
												.valid_out(per_bank_mem_rsp_valid),
												.data_out(per_bank_mem_rsp_pdata),
												.sel_out(),
												.ready_out(per_bank_mem_rsp_ready),
												.collisions()
											);
											// Trace: src/VX_cache.sv:146:5
											wire [511:0] per_bank_mem_rsp_data;
											// Trace: src/VX_cache.sv:147:5
											wire [4:0] per_bank_mem_rsp_tag;
											// Trace: src/VX_cache.sv:148:5
											genvar _gv_i_32;
											for (_gv_i_32 = 0; _gv_i_32 < NUM_BANKS; _gv_i_32 = _gv_i_32 + 1) begin : g_per_bank_mem_rsp_data
												localparam i = _gv_i_32;
												// Trace: src/VX_cache.sv:149:9
												assign {per_bank_mem_rsp_data[i * 512+:512], per_bank_mem_rsp_tag[i * 5+:5]} = per_bank_mem_rsp_pdata[i * 517+:517];
											end
											// Trace: src/VX_cache.sv:154:5
											wire [0:0] per_bank_core_req_valid;
											// Trace: src/VX_cache.sv:155:5
											wire [25:0] per_bank_core_req_addr;
											// Trace: src/VX_cache.sv:156:5
											wire [0:0] per_bank_core_req_rw;
											// Trace: src/VX_cache.sv:157:5
											wire [3:0] per_bank_core_req_wsel;
											// Trace: src/VX_cache.sv:158:5
											wire [3:0] per_bank_core_req_byteen;
											// Trace: src/VX_cache.sv:159:5
											wire [31:0] per_bank_core_req_data;
											// Trace: src/VX_cache.sv:160:5
											wire [2:0] per_bank_core_req_tag;
											// Trace: src/VX_cache.sv:161:5
											wire [0:0] per_bank_core_req_idx;
											// Trace: src/VX_cache.sv:162:5
											wire [0:0] per_bank_core_req_flags;
											// Trace: src/VX_cache.sv:163:5
											wire [0:0] per_bank_core_req_ready;
											// Trace: src/VX_cache.sv:164:5
											wire [0:0] per_bank_core_rsp_valid;
											// Trace: src/VX_cache.sv:165:5
											wire [31:0] per_bank_core_rsp_data;
											// Trace: src/VX_cache.sv:166:5
											wire [2:0] per_bank_core_rsp_tag;
											// Trace: src/VX_cache.sv:167:5
											wire [0:0] per_bank_core_rsp_idx;
											// Trace: src/VX_cache.sv:168:5
											wire [0:0] per_bank_core_rsp_ready;
											// Trace: src/VX_cache.sv:169:5
											wire [0:0] per_bank_mem_req_valid;
											// Trace: src/VX_cache.sv:170:5
											wire [25:0] per_bank_mem_req_addr;
											// Trace: src/VX_cache.sv:171:5
											wire [0:0] per_bank_mem_req_rw;
											// Trace: src/VX_cache.sv:172:5
											wire [63:0] per_bank_mem_req_byteen;
											// Trace: src/VX_cache.sv:173:5
											wire [511:0] per_bank_mem_req_data;
											// Trace: src/VX_cache.sv:174:5
											wire [4:0] per_bank_mem_req_tag;
											// Trace: src/VX_cache.sv:175:5
											wire [0:0] per_bank_mem_req_flags;
											// Trace: src/VX_cache.sv:176:5
											wire [0:0] per_bank_mem_req_ready;
											// Trace: src/VX_cache.sv:177:5
											wire [0:0] core_req_valid;
											// Trace: src/VX_cache.sv:178:5
											wire [29:0] core_req_addr;
											// Trace: src/VX_cache.sv:179:5
											wire [0:0] core_req_rw;
											// Trace: src/VX_cache.sv:180:5
											wire [3:0] core_req_byteen;
											// Trace: src/VX_cache.sv:181:5
											wire [31:0] core_req_data;
											// Trace: src/VX_cache.sv:182:5
											wire [2:0] core_req_tag;
											// Trace: src/VX_cache.sv:183:5
											wire [0:0] core_req_flags;
											// Trace: src/VX_cache.sv:184:5
											wire [0:0] core_req_ready;
											// Trace: src/VX_cache.sv:185:5
											wire [25:0] core_req_line_addr;
											// Trace: src/VX_cache.sv:186:5
											wire [0:0] core_req_bid;
											// Trace: src/VX_cache.sv:187:5
											wire [3:0] core_req_wsel;
											// Trace: src/VX_cache.sv:188:5
											wire [70:0] core_req_data_in;
											// Trace: src/VX_cache.sv:189:5
											wire [70:0] core_req_data_out;
											// Trace: src/VX_cache.sv:190:5
											genvar _gv_i_33;
											for (_gv_i_33 = 0; _gv_i_33 < NUM_REQS; _gv_i_33 = _gv_i_33 + 1) begin : g_core_req
												localparam i = _gv_i_33;
												// Trace: src/VX_cache.sv:191:9
												assign core_req_valid[i] = core_bus2_if[i].req_valid;
												// Trace: src/VX_cache.sv:192:9
												assign core_req_rw[i] = core_bus2_if[i].req_data[72];
												// Trace: src/VX_cache.sv:193:9
												assign core_req_byteen[i * 4+:4] = core_bus2_if[i].req_data[9-:4];
												// Trace: src/VX_cache.sv:194:9
												assign core_req_addr[i * 30+:30] = core_bus2_if[i].req_data[71-:30];
												// Trace: src/VX_cache.sv:195:9
												assign core_req_data[i * 32+:32] = core_bus2_if[i].req_data[41-:32];
												// Trace: src/VX_cache.sv:196:9
												assign core_req_tag[i * 3+:3] = core_bus2_if[i].req_data[2-:3];
												// Trace: src/VX_cache.sv:197:9
												assign core_req_flags[i+:1] = sv2v_cast_1(core_bus2_if[i].req_data[5-:3]);
												// Trace: src/VX_cache.sv:198:9
												assign core_bus2_if[i].req_ready = core_req_ready[i];
											end
											// Trace: src/VX_cache.sv:200:5
											genvar _gv_i_34;
											for (_gv_i_34 = 0; _gv_i_34 < NUM_REQS; _gv_i_34 = _gv_i_34 + 1) begin : g_core_req_wsel
												localparam i = _gv_i_34;
												if (1) begin : g_wsel
													// Trace: src/VX_cache.sv:202:13
													assign core_req_wsel[i * 4+:4] = core_req_addr[i * 30+:WORD_SEL_BITS];
												end
											end
											// Trace: src/VX_cache.sv:207:5
											genvar _gv_i_35;
											for (_gv_i_35 = 0; _gv_i_35 < NUM_REQS; _gv_i_35 = _gv_i_35 + 1) begin : g_core_req_line_addr
												localparam i = _gv_i_35;
												// Trace: src/VX_cache.sv:208:9
												assign core_req_line_addr[i * 26+:26] = core_req_addr[(i * 30) + 4+:LINE_ADDR_WIDTH];
											end
											// Trace: src/VX_cache.sv:210:5
											genvar _gv_i_36;
											for (_gv_i_36 = 0; _gv_i_36 < NUM_REQS; _gv_i_36 = _gv_i_36 + 1) begin : g_core_req_bid
												localparam i = _gv_i_36;
												if (1) begin : g_singlebank
													// Trace: src/VX_cache.sv:214:13
													assign core_req_bid[i+:1] = 1'sb0;
												end
											end
											// Trace: src/VX_cache.sv:217:5
											genvar _gv_i_37;
											for (_gv_i_37 = 0; _gv_i_37 < NUM_REQS; _gv_i_37 = _gv_i_37 + 1) begin : g_core_req_data_in
												localparam i = _gv_i_37;
												// Trace: src/VX_cache.sv:218:9
												assign core_req_data_in[i * 71+:71] = {core_req_line_addr[i * 26+:26], core_req_rw[i], core_req_wsel[i * 4+:4], core_req_byteen[i * 4+:4], core_req_data[i * 32+:32], core_req_tag[i * 3+:3], core_req_flags[i+:1]};
											end
											// Trace: src/VX_cache.sv:228:5
											assign per_bank_core_req_fire = per_bank_core_req_valid & per_bank_mem_req_ready;
											// Trace: src/VX_cache.sv:229:5
											VX_stream_xbar #(
												.NUM_INPUTS(NUM_REQS),
												.NUM_OUTPUTS(NUM_BANKS),
												.DATAW(CORE_REQ_DATAW),
												.PERF_CTR_BITS(44),
												.ARBITER("R"),
												.OUT_BUF(REQ_XBAR_BUF)
											) req_xbar(
												.clk(clk),
												.reset(reset),
												.collisions(),
												.valid_in(core_req_valid),
												.data_in(core_req_data_in),
												.sel_in(core_req_bid),
												.ready_in(core_req_ready),
												.valid_out(per_bank_core_req_valid),
												.data_out(core_req_data_out),
												.sel_out(per_bank_core_req_idx),
												.ready_out(per_bank_core_req_ready)
											);
											// Trace: src/VX_cache.sv:249:5
											genvar _gv_i_38;
											for (_gv_i_38 = 0; _gv_i_38 < NUM_BANKS; _gv_i_38 = _gv_i_38 + 1) begin : g_core_req_data_out
												localparam i = _gv_i_38;
												// Trace: src/VX_cache.sv:250:9
												assign {per_bank_core_req_addr[i * 26+:26], per_bank_core_req_rw[i], per_bank_core_req_wsel[i * 4+:4], per_bank_core_req_byteen[i * 4+:4], per_bank_core_req_data[i * 32+:32], per_bank_core_req_tag[i * 3+:3], per_bank_core_req_flags[i+:1]} = core_req_data_out[i * 71+:71];
											end
											// Trace: src/VX_cache.sv:260:5
											genvar _gv_bank_id_1;
											for (_gv_bank_id_1 = 0; _gv_bank_id_1 < NUM_BANKS; _gv_bank_id_1 = _gv_bank_id_1 + 1) begin : g_banks
												localparam bank_id = _gv_bank_id_1;
												// Trace: src/VX_cache.sv:261:9
												VX_cache_bank #(
													.BANK_ID(bank_id),
													.INSTANCE_ID(""),
													.CACHE_SIZE(CACHE_SIZE),
													.LINE_SIZE(LINE_SIZE),
													.NUM_BANKS(NUM_BANKS),
													.NUM_WAYS(NUM_WAYS),
													.WORD_SIZE(WORD_SIZE),
													.NUM_REQS(NUM_REQS),
													.WRITE_ENABLE(WRITE_ENABLE),
													.WRITEBACK(WRITEBACK),
													.DIRTY_BYTES(DIRTY_BYTES),
													.REPL_POLICY(REPL_POLICY),
													.CRSQ_SIZE(CRSQ_SIZE),
													.MSHR_SIZE(MSHR_SIZE),
													.MREQ_SIZE(MREQ_SIZE),
													.UUID_WIDTH(UUID_WIDTH),
													.TAG_WIDTH(TAG_WIDTH),
													.FLAGS_WIDTH(FLAGS_WIDTH),
													.CORE_OUT_REG((CORE_RSP_REG_DISABLE ? 0 : 1)),
													.MEM_OUT_REG((MEM_REQ_REG_DISABLE ? 0 : 1))
												) bank(
													.clk(clk),
													.reset(reset),
													.core_req_valid(per_bank_core_req_valid[bank_id]),
													.core_req_addr(per_bank_core_req_addr[bank_id * 26+:26]),
													.core_req_rw(per_bank_core_req_rw[bank_id]),
													.core_req_wsel(per_bank_core_req_wsel[bank_id * 4+:4]),
													.core_req_byteen(per_bank_core_req_byteen[bank_id * 4+:4]),
													.core_req_data(per_bank_core_req_data[bank_id * 32+:32]),
													.core_req_tag(per_bank_core_req_tag[bank_id * 3+:3]),
													.core_req_idx(per_bank_core_req_idx[bank_id+:1]),
													.core_req_flags(per_bank_core_req_flags[bank_id+:1]),
													.core_req_ready(per_bank_core_req_ready[bank_id]),
													.core_rsp_valid(per_bank_core_rsp_valid[bank_id]),
													.core_rsp_data(per_bank_core_rsp_data[bank_id * 32+:32]),
													.core_rsp_tag(per_bank_core_rsp_tag[bank_id * 3+:3]),
													.core_rsp_idx(per_bank_core_rsp_idx[bank_id+:1]),
													.core_rsp_ready(per_bank_core_rsp_ready[bank_id]),
													.mem_req_valid(per_bank_mem_req_valid[bank_id]),
													.mem_req_addr(per_bank_mem_req_addr[bank_id * 26+:26]),
													.mem_req_rw(per_bank_mem_req_rw[bank_id]),
													.mem_req_byteen(per_bank_mem_req_byteen[bank_id * 64+:64]),
													.mem_req_data(per_bank_mem_req_data[bank_id * 512+:512]),
													.mem_req_tag(per_bank_mem_req_tag[bank_id * 5+:5]),
													.mem_req_flags(per_bank_mem_req_flags[bank_id+:1]),
													.mem_req_ready(per_bank_mem_req_ready[bank_id]),
													.mem_rsp_valid(per_bank_mem_rsp_valid[bank_id]),
													.mem_rsp_data(per_bank_mem_rsp_data[bank_id * 512+:512]),
													.mem_rsp_tag(per_bank_mem_rsp_tag[bank_id * 5+:5]),
													.mem_rsp_ready(per_bank_mem_rsp_ready[bank_id]),
													.flush_begin(per_bank_flush_begin[bank_id]),
													.flush_uuid(flush_uuid),
													.flush_end(per_bank_flush_end[bank_id])
												);
											end
											// Trace: src/VX_cache.sv:317:5
											wire [34:0] core_rsp_data_in;
											// Trace: src/VX_cache.sv:318:5
											wire [34:0] core_rsp_data_out;
											// Trace: src/VX_cache.sv:319:5
											wire [0:0] core_rsp_valid_s;
											// Trace: src/VX_cache.sv:320:5
											wire [31:0] core_rsp_data_s;
											// Trace: src/VX_cache.sv:321:5
											wire [2:0] core_rsp_tag_s;
											// Trace: src/VX_cache.sv:322:5
											wire [0:0] core_rsp_ready_s;
											// Trace: src/VX_cache.sv:323:5
											genvar _gv_i_39;
											for (_gv_i_39 = 0; _gv_i_39 < NUM_BANKS; _gv_i_39 = _gv_i_39 + 1) begin : g_core_rsp_data_in
												localparam i = _gv_i_39;
												// Trace: src/VX_cache.sv:324:9
												assign core_rsp_data_in[i * 35+:35] = {per_bank_core_rsp_data[i * 32+:32], per_bank_core_rsp_tag[i * 3+:3]};
											end
											// Trace: src/VX_cache.sv:326:5
											VX_stream_xbar #(
												.NUM_INPUTS(NUM_BANKS),
												.NUM_OUTPUTS(NUM_REQS),
												.DATAW(CORE_RSP_DATAW),
												.ARBITER("R")
											) rsp_xbar(
												.clk(clk),
												.reset(reset),
												.collisions(),
												.valid_in(per_bank_core_rsp_valid),
												.data_in(core_rsp_data_in),
												.sel_in(per_bank_core_rsp_idx),
												.ready_in(per_bank_core_rsp_ready),
												.valid_out(core_rsp_valid_s),
												.data_out(core_rsp_data_out),
												.ready_out(core_rsp_ready_s),
												.sel_out()
											);
											// Trace: src/VX_cache.sv:344:5
											genvar _gv_i_40;
											for (_gv_i_40 = 0; _gv_i_40 < NUM_REQS; _gv_i_40 = _gv_i_40 + 1) begin : g_core_rsp_data_s
												localparam i = _gv_i_40;
												// Trace: src/VX_cache.sv:345:9
												assign {core_rsp_data_s[i * 32+:32], core_rsp_tag_s[i * 3+:3]} = core_rsp_data_out[i * 35+:35];
											end
											// Trace: src/VX_cache.sv:347:5
											genvar _gv_i_41;
											for (_gv_i_41 = 0; _gv_i_41 < NUM_REQS; _gv_i_41 = _gv_i_41 + 1) begin : g_core_rsp_buf
												localparam i = _gv_i_41;
												// Trace: src/VX_cache.sv:348:9
												VX_elastic_buffer #(
													.DATAW(35),
													.SIZE((CORE_RSP_REG_DISABLE ? ((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : 2) : 0)),
													.OUT_REG(((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : (CORE_OUT_BUF & 7) - 2))
												) core_rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(core_rsp_valid_s[i]),
													.ready_in(core_rsp_ready_s[i]),
													.data_in({core_rsp_data_s[i * 32+:32], core_rsp_tag_s[i * 3+:3]}),
													.data_out({core_bus2_if[i].rsp_data[34-:32], core_bus2_if[i].rsp_data[2-:3]}),
													.valid_out(core_bus2_if[i].rsp_valid),
													.ready_out(core_bus2_if[i].rsp_ready)
												);
											end
											// Trace: src/VX_cache.sv:363:5
											wire [608:0] per_bank_mem_req_pdata;
											// Trace: src/VX_cache.sv:364:5
											genvar _gv_i_42;
											for (_gv_i_42 = 0; _gv_i_42 < NUM_BANKS; _gv_i_42 = _gv_i_42 + 1) begin : g_per_bank_mem_req_pdata
												localparam i = _gv_i_42;
												// Trace: src/VX_cache.sv:365:9
												assign per_bank_mem_req_pdata[i * 609+:609] = {per_bank_mem_req_rw[i], per_bank_mem_req_addr[i * 26+:26], per_bank_mem_req_data[i * 512+:512], per_bank_mem_req_byteen[i * 64+:64], per_bank_mem_req_flags[i+:1], per_bank_mem_req_tag[i * 5+:5]};
											end
											// Trace: src/VX_cache.sv:374:5
											wire [0:0] mem_req_valid;
											// Trace: src/VX_cache.sv:375:5
											wire [608:0] mem_req_pdata;
											// Trace: src/VX_cache.sv:376:5
											wire [0:0] mem_req_ready;
											// Trace: src/VX_cache.sv:377:5
											wire [0:0] mem_req_sel_out;
											// Trace: src/VX_cache.sv:378:5
											VX_stream_arb #(
												.NUM_INPUTS(NUM_BANKS),
												.NUM_OUTPUTS(MEM_PORTS),
												.DATAW(MEM_REQ_DATAW),
												.ARBITER("R")
											) mem_req_arb(
												.clk(clk),
												.reset(reset),
												.valid_in(per_bank_mem_req_valid),
												.data_in(per_bank_mem_req_pdata),
												.ready_in(per_bank_mem_req_ready),
												.valid_out(mem_req_valid),
												.data_out(mem_req_pdata),
												.ready_out(mem_req_ready),
												.sel_out(mem_req_sel_out)
											);
											// Trace: src/VX_cache.sv:394:5
											genvar _gv_i_43;
											for (_gv_i_43 = 0; _gv_i_43 < MEM_PORTS; _gv_i_43 = _gv_i_43 + 1) begin : g_mem_req_buf
												localparam i = _gv_i_43;
												// Trace: src/VX_cache.sv:395:9
												wire mem_req_rw;
												// Trace: src/VX_cache.sv:396:9
												wire [25:0] mem_req_addr;
												// Trace: src/VX_cache.sv:397:9
												wire [511:0] mem_req_data;
												// Trace: src/VX_cache.sv:398:9
												wire [63:0] mem_req_byteen;
												// Trace: src/VX_cache.sv:399:9
												wire [0:0] mem_req_flags;
												// Trace: src/VX_cache.sv:400:9
												wire [4:0] mem_req_tag;
												// Trace: src/VX_cache.sv:401:9
												assign {mem_req_rw, mem_req_addr, mem_req_data, mem_req_byteen, mem_req_flags, mem_req_tag} = mem_req_pdata[i * 609+:609];
												// Trace: src/VX_cache.sv:409:9
												wire [25:0] mem_req_addr_w;
												// Trace: src/VX_cache.sv:410:9
												wire [4:0] mem_req_tag_w;
												// Trace: src/VX_cache.sv:411:9
												wire [0:0] mem_req_flags_w;
												if (1) begin : g_mem_req_tag
													// Trace: src/VX_cache.sv:430:13
													assign mem_req_addr_w = mem_req_addr;
													// Trace: src/VX_cache.sv:431:13
													assign mem_req_tag_w = mem_req_tag;
												end
												// Trace: src/VX_cache.sv:433:9
												VX_elastic_buffer #(
													.DATAW(609),
													.SIZE((MEM_REQ_REG_DISABLE ? ((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : 2) : 0)),
													.OUT_REG(((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : (MEM_OUT_BUF & 7) - 2))
												) mem_req_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_req_valid[i]),
													.ready_in(mem_req_ready[i]),
													.data_in({mem_req_rw, mem_req_byteen, mem_req_addr_w, mem_req_data, mem_req_tag_w, mem_req_flags}),
													.data_out({mem_bus_tmp_if[i].req_data[610], mem_bus_tmp_if[i].req_data[71-:64], mem_bus_tmp_if[i].req_data[609-:26], mem_bus_tmp_if[i].req_data[583-:512], mem_bus_tmp_if[i].req_data[4-:5], mem_req_flags_w}),
													.valid_out(mem_bus_tmp_if[i].req_valid),
													.ready_out(mem_bus_tmp_if[i].req_ready)
												);
												if (1) begin : g_no_mem_req_flags
													// Trace: src/VX_cache.sv:450:13
													assign mem_bus_tmp_if[i].req_data[7-:3] = 1'sb0;
												end
												if (WRITE_ENABLE) begin : g_mem_bus_if
													// Trace: src/VX_cache.sv:453:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
													// Trace: src/VX_cache.sv:454:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
													// Trace: src/VX_cache.sv:455:5
													assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_ready;
													// Trace: src/VX_cache.sv:456:5
													assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_valid;
													// Trace: src/VX_cache.sv:457:5
													assign mem_bus_tmp_if[i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data;
													// Trace: src/VX_cache.sv:458:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
												end
												else begin : g_mem_bus_if_ro
													// Trace: src/VX_cache.sv:460:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
													// Trace: src/VX_cache.sv:461:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[610] = 0;
													// Trace: src/VX_cache.sv:462:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[609-:26] = mem_bus_tmp_if[i].req_data[609-:26];
													// Trace: src/VX_cache.sv:463:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[583-:512] = 1'sb0;
													// Trace: src/VX_cache.sv:464:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[71-:64] = 1'sb1;
													// Trace: src/VX_cache.sv:465:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[7-:3] = mem_bus_tmp_if[i].req_data[7-:3];
													// Trace: src/VX_cache.sv:466:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[4-:5] = mem_bus_tmp_if[i].req_data[4-:5];
													// Trace: src/VX_cache.sv:467:5
													assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_ready;
													// Trace: src/VX_cache.sv:468:5
													assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_valid;
													// Trace: src/VX_cache.sv:469:5
													assign mem_bus_tmp_if[i].rsp_data[516-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data[516-:512];
													// Trace: src/VX_cache.sv:470:5
													assign mem_bus_tmp_if[i].rsp_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data[4-:5];
													// Trace: src/VX_cache.sv:471:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
												end
											end
										end
										assign cache.clk = clk;
										assign cache.reset = reset;
									end
								end
								assign cache_wrap.clk = clk;
								assign cache_wrap.reset = reset;
							end
							// Trace: src/VX_cache_cluster.sv:124:5
							genvar _gv_i_67;
							for (_gv_i_67 = 0; _gv_i_67 < MEM_PORTS; _gv_i_67 = _gv_i_67 + 1) begin : g_mem_bus_if
								localparam i = _gv_i_67;
								// Trace: src/VX_cache_cluster.sv:125:9
								// expanded interface instance: arb_core_bus_tmp_if
								localparam _param_E788B_DATA_SIZE = LINE_SIZE;
								localparam _param_E788B_TAG_WIDTH = MEM_TAG_WIDTH;
								genvar _arr_E788B;
								for (_arr_E788B = 0; _arr_E788B <= 0; _arr_E788B = _arr_E788B + 1) begin : arb_core_bus_tmp_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_E788B_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_E788B_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [610:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [516:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								// Trace: src/VX_cache_cluster.sv:129:9
								// expanded interface instance: mem_bus_tmp_if
								localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
								localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH + 0;
								genvar _arr_4FE36;
								for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [610:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [516:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								genvar _gv_j_7;
								for (_gv_j_7 = 0; _gv_j_7 < NUM_CACHES; _gv_j_7 = _gv_j_7 + 1) begin : g_arb_core_bus_tmp_if
									localparam j = _gv_j_7;
									// Trace: src/VX_cache_cluster.sv:134:5
									assign arb_core_bus_tmp_if[j].req_valid = cache_mem_bus_if[(j * MEM_PORTS) + i].req_valid;
									// Trace: src/VX_cache_cluster.sv:135:5
									assign arb_core_bus_tmp_if[j].req_data = cache_mem_bus_if[(j * MEM_PORTS) + i].req_data;
									// Trace: src/VX_cache_cluster.sv:136:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].req_ready = arb_core_bus_tmp_if[j].req_ready;
									// Trace: src/VX_cache_cluster.sv:137:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_valid = arb_core_bus_tmp_if[j].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:138:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_data = arb_core_bus_tmp_if[j].rsp_data;
									// Trace: src/VX_cache_cluster.sv:139:5
									assign arb_core_bus_tmp_if[j].rsp_ready = cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_ready;
								end
								// Trace: src/VX_cache_cluster.sv:141:9
								// expanded module instance: mem_arb
								localparam _bbase_7277A_bus_in_if = 0;
								localparam _bbase_7277A_bus_out_if = 0;
								localparam _param_7277A_NUM_INPUTS = NUM_CACHES;
								localparam _param_7277A_NUM_OUTPUTS = 1;
								localparam _param_7277A_DATA_SIZE = LINE_SIZE;
								localparam _param_7277A_TAG_WIDTH = MEM_TAG_WIDTH;
								localparam _param_7277A_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_7277A_ARBITER = "R";
								localparam _param_7277A_REQ_OUT_BUF = 0;
								localparam _param_7277A_RSP_OUT_BUF = 0;
								if (1) begin : mem_arb
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_7277A_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = _param_7277A_NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_7277A_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_7277A_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_7277A_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_7277A_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_7277A_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:16
									localparam ARBITER = _param_7277A_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 512;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 0;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 606 + TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [0:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [REQ_DATAW - 1:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [0:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [REQ_DATAW - 1:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_80;
									for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
										localparam i = _gv_i_80;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 611+:611] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_81;
									for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
										localparam i = _gv_i_81;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [TAG_WIDTH - 1:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										VX_bits_insert #(
											.N(TAG_WIDTH),
											.S(LOG_NUM_REQS),
											.POS(TAG_SEL_IDX)
										) bits_insert(
											.data_in(req_tag_out),
											.ins_in(req_sel_out[i+:1]),
											.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[4-:5])
										);
										// Trace: src/VX_mem_arb.sv:64:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:65:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[610], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[609-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[583-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[71-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[7-:3], req_tag_out} = req_data_out[i * 611+:611];
										// Trace: src/VX_mem_arb.sv:73:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
									end
									// Trace: src/VX_mem_arb.sv:75:5
									wire [0:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:76:5
									wire [RSP_DATAW - 1:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:77:5
									wire [0:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:78:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:79:5
									wire [RSP_DATAW - 1:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:81:5
									if (1) begin : g_passthru
										genvar _gv_i_83;
										for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_83;
											// Trace: src/VX_mem_arb.sv:116:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:117:13
											assign rsp_data_in[i * 517+:517] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
											// Trace: src/VX_mem_arb.sv:118:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:120:9
										VX_stream_arb #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.ARBITER(ARBITER),
											.OUT_BUF(RSP_OUT_BUF)
										) req_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
									end
									// Trace: src/VX_mem_arb.sv:138:5
									genvar _gv_i_84;
									for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
										localparam i = _gv_i_84;
										// Trace: src/VX_mem_arb.sv:139:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:140:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 517+:517];
										// Trace: src/VX_mem_arb.sv:141:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign mem_arb.clk = clk;
								assign mem_arb.reset = reset;
								if (WRITE_ENABLE) begin : g_we
									// Trace: src/VX_cache_cluster.sv:157:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[0].req_valid;
									// Trace: src/VX_cache_cluster.sv:158:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[0].req_data;
									// Trace: src/VX_cache_cluster.sv:159:5
									assign mem_bus_tmp_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
									// Trace: src/VX_cache_cluster.sv:160:5
									assign mem_bus_tmp_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:161:5
									assign mem_bus_tmp_if[0].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
									// Trace: src/VX_cache_cluster.sv:162:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[0].rsp_ready;
								end
								else begin : g_ro
									// Trace: src/VX_cache_cluster.sv:164:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[0].req_valid;
									// Trace: src/VX_cache_cluster.sv:165:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[610] = 0;
									// Trace: src/VX_cache_cluster.sv:166:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[609-:26] = mem_bus_tmp_if[0].req_data[609-:26];
									// Trace: src/VX_cache_cluster.sv:167:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[583-:512] = 1'sb0;
									// Trace: src/VX_cache_cluster.sv:168:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[71-:64] = 1'sb1;
									// Trace: src/VX_cache_cluster.sv:169:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[7-:3] = mem_bus_tmp_if[0].req_data[7-:3];
									// Trace: src/VX_cache_cluster.sv:170:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[4-:5] = mem_bus_tmp_if[0].req_data[4-:5];
									// Trace: src/VX_cache_cluster.sv:171:5
									assign mem_bus_tmp_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
									// Trace: src/VX_cache_cluster.sv:172:5
									assign mem_bus_tmp_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:173:5
									assign mem_bus_tmp_if[0].rsp_data[516-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[516-:512];
									// Trace: src/VX_cache_cluster.sv:174:5
									assign mem_bus_tmp_if[0].rsp_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[4-:5];
									// Trace: src/VX_cache_cluster.sv:175:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[0].rsp_ready;
								end
							end
						end
						assign icache.clk = clk;
						assign icache.reset = icache_reset;
						// Trace: src/VX_socket.sv:55:5
						localparam VX_gpu_pkg_DCACHE_MERGED_REQS = 1;
						localparam VX_gpu_pkg_DCACHE_MEM_BATCHES = 1;
						localparam VX_gpu_pkg_DCACHE_TAG_ID_BITS = 2;
						localparam VX_gpu_pkg_DCACHE_TAG_WIDTH = 3;
						// expanded interface instance: per_core_dcache_bus_if
						localparam _param_F6DD5_DATA_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
						localparam _param_F6DD5_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
						genvar _arr_F6DD5;
						for (_arr_F6DD5 = 0; _arr_F6DD5 <= 0; _arr_F6DD5 = _arr_F6DD5 + 1) begin : per_core_dcache_bus_if
							// Trace: src/VX_mem_bus_if.sv:2:15
							localparam DATA_SIZE = _param_F6DD5_DATA_SIZE;
							// Trace: src/VX_mem_bus_if.sv:3:15
							localparam FLAGS_WIDTH = 3;
							// Trace: src/VX_mem_bus_if.sv:4:15
							localparam TAG_WIDTH = _param_F6DD5_TAG_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:5:15
							localparam MEM_ADDR_WIDTH = 32;
							// Trace: src/VX_mem_bus_if.sv:6:15
							localparam ADDR_WIDTH = 28;
							// Trace: src/VX_mem_bus_if.sv:7:15
							localparam UUID_WIDTH = 1;
							// Trace: src/VX_mem_bus_if.sv:9:5
							// removed localparam type tag_t
							// Trace: src/VX_mem_bus_if.sv:13:5
							// removed localparam type req_data_t
							// Trace: src/VX_mem_bus_if.sv:21:5
							// removed localparam type rsp_data_t
							// Trace: src/VX_mem_bus_if.sv:25:5
							wire req_valid;
							// Trace: src/VX_mem_bus_if.sv:26:5
							wire [178:0] req_data;
							// Trace: src/VX_mem_bus_if.sv:27:5
							wire req_ready;
							// Trace: src/VX_mem_bus_if.sv:28:5
							wire rsp_valid;
							// Trace: src/VX_mem_bus_if.sv:29:5
							wire [130:0] rsp_data;
							// Trace: src/VX_mem_bus_if.sv:30:5
							wire rsp_ready;
							// Trace: src/VX_mem_bus_if.sv:31:5
							// Trace: src/VX_mem_bus_if.sv:39:5
						end
						// Trace: src/VX_socket.sv:59:5
						localparam VX_gpu_pkg_DCACHE_LINE_SIZE = 64;
						localparam VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH = 6;
						// expanded interface instance: dcache_mem_bus_if
						localparam _param_28DB2_DATA_SIZE = VX_gpu_pkg_DCACHE_LINE_SIZE;
						localparam _param_28DB2_TAG_WIDTH = VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH;
						genvar _arr_28DB2;
						for (_arr_28DB2 = 0; _arr_28DB2 <= 0; _arr_28DB2 = _arr_28DB2 + 1) begin : dcache_mem_bus_if
							// Trace: src/VX_mem_bus_if.sv:2:15
							localparam DATA_SIZE = _param_28DB2_DATA_SIZE;
							// Trace: src/VX_mem_bus_if.sv:3:15
							localparam FLAGS_WIDTH = 3;
							// Trace: src/VX_mem_bus_if.sv:4:15
							localparam TAG_WIDTH = _param_28DB2_TAG_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:5:15
							localparam MEM_ADDR_WIDTH = 32;
							// Trace: src/VX_mem_bus_if.sv:6:15
							localparam ADDR_WIDTH = 26;
							// Trace: src/VX_mem_bus_if.sv:7:15
							localparam UUID_WIDTH = 1;
							// Trace: src/VX_mem_bus_if.sv:9:5
							// removed localparam type tag_t
							// Trace: src/VX_mem_bus_if.sv:13:5
							// removed localparam type req_data_t
							// Trace: src/VX_mem_bus_if.sv:21:5
							// removed localparam type rsp_data_t
							// Trace: src/VX_mem_bus_if.sv:25:5
							wire req_valid;
							// Trace: src/VX_mem_bus_if.sv:26:5
							wire [611:0] req_data;
							// Trace: src/VX_mem_bus_if.sv:27:5
							wire req_ready;
							// Trace: src/VX_mem_bus_if.sv:28:5
							wire rsp_valid;
							// Trace: src/VX_mem_bus_if.sv:29:5
							wire [517:0] rsp_data;
							// Trace: src/VX_mem_bus_if.sv:30:5
							wire rsp_ready;
							// Trace: src/VX_mem_bus_if.sv:31:5
							// Trace: src/VX_mem_bus_if.sv:39:5
						end
						// Trace: src/VX_socket.sv:63:5
						wire [0:0] dcache_reset;
						// Trace: src/VX_socket.sv:64:5
						VX_reset_relay #(
							.N(1),
							.MAX_FANOUT(0)
						) __dcache_reset(
							.clk(clk),
							.reset(reset),
							.reset_o(dcache_reset)
						);
						// Trace: src/VX_socket.sv:69:5
						// expanded module instance: dcache
						localparam _bbase_CC492_core_bus_if = 0;
						localparam _bbase_CC492_mem_bus_if = 0;
						localparam _param_CC492_INSTANCE_ID = "";
						localparam _param_CC492_NUM_UNITS = 1;
						localparam _param_CC492_NUM_INPUTS = 1;
						localparam _param_CC492_TAG_SEL_IDX = 0;
						localparam _param_CC492_CACHE_SIZE = 16384;
						localparam _param_CC492_LINE_SIZE = VX_gpu_pkg_DCACHE_LINE_SIZE;
						localparam _param_CC492_NUM_BANKS = VX_gpu_pkg_DCACHE_NUM_REQS;
						localparam _param_CC492_NUM_WAYS = 4;
						localparam _param_CC492_WORD_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
						localparam _param_CC492_NUM_REQS = VX_gpu_pkg_DCACHE_NUM_REQS;
						localparam _param_CC492_MEM_PORTS = VX_gpu_pkg_DCACHE_NUM_REQS;
						localparam _param_CC492_CRSQ_SIZE = 2;
						localparam _param_CC492_MSHR_SIZE = 16;
						localparam _param_CC492_MRSQ_SIZE = 4;
						localparam _param_CC492_MREQ_SIZE = 4;
						localparam _param_CC492_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
						localparam _param_CC492_UUID_WIDTH = 1;
						localparam _param_CC492_FLAGS_WIDTH = 3;
						localparam _param_CC492_WRITE_ENABLE = 1;
						localparam _param_CC492_WRITEBACK = 0;
						localparam _param_CC492_DIRTY_BYTES = 0;
						localparam _param_CC492_REPL_POLICY = 1;
						localparam _param_CC492_NC_ENABLE = 1;
						localparam _param_CC492_CORE_OUT_BUF = 3;
						localparam _param_CC492_MEM_OUT_BUF = 2;
						if (1) begin : dcache
							// removed import VX_gpu_pkg::*;
							// Trace: src/VX_cache_cluster.sv:2:16
							localparam INSTANCE_ID = _param_CC492_INSTANCE_ID;
							// Trace: src/VX_cache_cluster.sv:3:15
							localparam NUM_UNITS = _param_CC492_NUM_UNITS;
							// Trace: src/VX_cache_cluster.sv:4:15
							localparam NUM_INPUTS = _param_CC492_NUM_INPUTS;
							// Trace: src/VX_cache_cluster.sv:5:15
							localparam TAG_SEL_IDX = _param_CC492_TAG_SEL_IDX;
							// Trace: src/VX_cache_cluster.sv:6:15
							localparam NUM_REQS = _param_CC492_NUM_REQS;
							// Trace: src/VX_cache_cluster.sv:7:15
							localparam MEM_PORTS = _param_CC492_MEM_PORTS;
							// Trace: src/VX_cache_cluster.sv:8:15
							localparam CACHE_SIZE = _param_CC492_CACHE_SIZE;
							// Trace: src/VX_cache_cluster.sv:9:15
							localparam LINE_SIZE = _param_CC492_LINE_SIZE;
							// Trace: src/VX_cache_cluster.sv:10:15
							localparam NUM_BANKS = _param_CC492_NUM_BANKS;
							// Trace: src/VX_cache_cluster.sv:11:15
							localparam NUM_WAYS = _param_CC492_NUM_WAYS;
							// Trace: src/VX_cache_cluster.sv:12:15
							localparam WORD_SIZE = _param_CC492_WORD_SIZE;
							// Trace: src/VX_cache_cluster.sv:13:15
							localparam CRSQ_SIZE = _param_CC492_CRSQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:14:15
							localparam MSHR_SIZE = _param_CC492_MSHR_SIZE;
							// Trace: src/VX_cache_cluster.sv:15:15
							localparam MRSQ_SIZE = _param_CC492_MRSQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:16:15
							localparam MREQ_SIZE = _param_CC492_MREQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:17:15
							localparam WRITE_ENABLE = _param_CC492_WRITE_ENABLE;
							// Trace: src/VX_cache_cluster.sv:18:15
							localparam WRITEBACK = _param_CC492_WRITEBACK;
							// Trace: src/VX_cache_cluster.sv:19:15
							localparam DIRTY_BYTES = _param_CC492_DIRTY_BYTES;
							// Trace: src/VX_cache_cluster.sv:20:15
							localparam REPL_POLICY = _param_CC492_REPL_POLICY;
							// Trace: src/VX_cache_cluster.sv:21:15
							localparam UUID_WIDTH = _param_CC492_UUID_WIDTH;
							// Trace: src/VX_cache_cluster.sv:22:15
							localparam TAG_WIDTH = _param_CC492_TAG_WIDTH;
							// Trace: src/VX_cache_cluster.sv:23:15
							localparam FLAGS_WIDTH = _param_CC492_FLAGS_WIDTH;
							// Trace: src/VX_cache_cluster.sv:24:15
							localparam NC_ENABLE = _param_CC492_NC_ENABLE;
							// Trace: src/VX_cache_cluster.sv:25:15
							localparam CORE_OUT_BUF = _param_CC492_CORE_OUT_BUF;
							// Trace: src/VX_cache_cluster.sv:26:15
							localparam MEM_OUT_BUF = _param_CC492_MEM_OUT_BUF;
							// Trace: src/VX_cache_cluster.sv:28:5
							wire clk;
							// Trace: src/VX_cache_cluster.sv:29:5
							wire reset;
							// Trace: src/VX_cache_cluster.sv:30:5
							localparam _mbase_core_bus_if = 0;
							// Trace: src/VX_cache_cluster.sv:31:5
							localparam _mbase_mem_bus_if = 0;
							// Trace: src/VX_cache_cluster.sv:33:5
							localparam NUM_CACHES = NUM_UNITS;
							// Trace: src/VX_cache_cluster.sv:34:5
							localparam PASSTHRU = 1'd0;
							// Trace: src/VX_cache_cluster.sv:35:5
							localparam ARB_TAG_WIDTH = 3;
							// Trace: src/VX_cache_cluster.sv:36:5
							localparam CACHE_MEM_TAG_WIDTH = 5;
							// Trace: src/VX_cache_cluster.sv:38:5
							localparam BYPASS_TAG_WIDTH = 5;
							// Trace: src/VX_cache_cluster.sv:40:5
							localparam NC_TAG_WIDTH = 6;
							// Trace: src/VX_cache_cluster.sv:41:5
							localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
							// Trace: src/VX_cache_cluster.sv:42:5
							// expanded interface instance: cache_mem_bus_if
							localparam _param_A4879_DATA_SIZE = LINE_SIZE;
							localparam _param_A4879_TAG_WIDTH = MEM_TAG_WIDTH;
							genvar _arr_A4879;
							for (_arr_A4879 = 0; _arr_A4879 <= 0; _arr_A4879 = _arr_A4879 + 1) begin : cache_mem_bus_if
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_A4879_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_A4879_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:7:15
								localparam UUID_WIDTH = 1;
								// Trace: src/VX_mem_bus_if.sv:9:5
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:13:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:21:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire [611:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire [517:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:30:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:31:5
								// Trace: src/VX_mem_bus_if.sv:39:5
							end
							// Trace: src/VX_cache_cluster.sv:46:5
							// expanded interface instance: arb_core_bus_if
							localparam _param_F9BC9_DATA_SIZE = WORD_SIZE;
							localparam _param_F9BC9_TAG_WIDTH = ARB_TAG_WIDTH;
							genvar _arr_F9BC9;
							for (_arr_F9BC9 = 0; _arr_F9BC9 <= 0; _arr_F9BC9 = _arr_F9BC9 + 1) begin : arb_core_bus_if
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_F9BC9_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam FLAGS_WIDTH = 3;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_F9BC9_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 28;
								// Trace: src/VX_mem_bus_if.sv:7:15
								localparam UUID_WIDTH = 1;
								// Trace: src/VX_mem_bus_if.sv:9:5
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:13:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:21:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire [178:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire [130:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:30:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:31:5
								// Trace: src/VX_mem_bus_if.sv:39:5
							end
							// Trace: src/VX_cache_cluster.sv:50:5
							genvar _gv_i_65;
							for (_gv_i_65 = 0; _gv_i_65 < NUM_REQS; _gv_i_65 = _gv_i_65 + 1) begin : g_core_arb
								localparam i = _gv_i_65;
								// Trace: src/VX_cache_cluster.sv:51:9
								// expanded interface instance: core_bus_tmp_if
								localparam _param_A62F7_DATA_SIZE = WORD_SIZE;
								localparam _param_A62F7_TAG_WIDTH = TAG_WIDTH;
								genvar _arr_A62F7;
								for (_arr_A62F7 = 0; _arr_A62F7 <= 0; _arr_A62F7 = _arr_A62F7 + 1) begin : core_bus_tmp_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_A62F7_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_A62F7_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 28;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [178:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [130:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								// Trace: src/VX_cache_cluster.sv:55:9
								// expanded interface instance: arb_core_bus_tmp_if
								localparam _param_E788B_DATA_SIZE = WORD_SIZE;
								localparam _param_E788B_TAG_WIDTH = ARB_TAG_WIDTH;
								genvar _arr_E788B;
								for (_arr_E788B = 0; _arr_E788B <= 0; _arr_E788B = _arr_E788B + 1) begin : arb_core_bus_tmp_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_E788B_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_E788B_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 28;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [178:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [130:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								genvar _gv_j_6;
								for (_gv_j_6 = 0; _gv_j_6 < NUM_INPUTS; _gv_j_6 = _gv_j_6 + 1) begin : g_core_bus_tmp_if
									localparam j = _gv_j_6;
									// Trace: src/VX_cache_cluster.sv:60:5
									assign core_bus_tmp_if[j].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_valid;
									// Trace: src/VX_cache_cluster.sv:61:5
									assign core_bus_tmp_if[j].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_data;
									// Trace: src/VX_cache_cluster.sv:62:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_ready = core_bus_tmp_if[j].req_ready;
									// Trace: src/VX_cache_cluster.sv:63:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_valid = core_bus_tmp_if[j].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:64:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_data = core_bus_tmp_if[j].rsp_data;
									// Trace: src/VX_cache_cluster.sv:65:5
									assign core_bus_tmp_if[j].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_ready;
								end
								// Trace: src/VX_cache_cluster.sv:67:9
								// expanded module instance: core_arb
								localparam _bbase_856A9_bus_in_if = 0;
								localparam _bbase_856A9_bus_out_if = 0;
								localparam _param_856A9_NUM_INPUTS = NUM_INPUTS;
								localparam _param_856A9_NUM_OUTPUTS = NUM_CACHES;
								localparam _param_856A9_DATA_SIZE = WORD_SIZE;
								localparam _param_856A9_TAG_WIDTH = TAG_WIDTH;
								localparam _param_856A9_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_856A9_ARBITER = "R";
								localparam _param_856A9_REQ_OUT_BUF = 0;
								localparam _param_856A9_RSP_OUT_BUF = 0;
								if (1) begin : core_arb
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_856A9_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = _param_856A9_NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_856A9_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_856A9_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_856A9_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_856A9_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_856A9_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:16
									localparam ARBITER = _param_856A9_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 28;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 128;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 0;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 179;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = 131;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [0:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [178:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [0:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [178:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_80;
									for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
										localparam i = _gv_i_80;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 179+:179] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_81;
									for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
										localparam i = _gv_i_81;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [2:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										VX_bits_insert #(
											.N(TAG_WIDTH),
											.S(LOG_NUM_REQS),
											.POS(TAG_SEL_IDX)
										) bits_insert(
											.data_in(req_tag_out),
											.ins_in(req_sel_out[i+:1]),
											.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[2-:3])
										);
										// Trace: src/VX_mem_arb.sv:64:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:65:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[178], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[177-:28], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[149-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[21-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[5-:3], req_tag_out} = req_data_out[i * 179+:179];
										// Trace: src/VX_mem_arb.sv:73:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
									end
									// Trace: src/VX_mem_arb.sv:75:5
									wire [0:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:76:5
									wire [130:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:77:5
									wire [0:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:78:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:79:5
									wire [130:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:81:5
									if (1) begin : g_passthru
										genvar _gv_i_83;
										for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_83;
											// Trace: src/VX_mem_arb.sv:116:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:117:13
											assign rsp_data_in[i * 131+:131] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
											// Trace: src/VX_mem_arb.sv:118:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:120:9
										VX_stream_arb #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.ARBITER(ARBITER),
											.OUT_BUF(RSP_OUT_BUF)
										) req_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
									end
									// Trace: src/VX_mem_arb.sv:138:5
									genvar _gv_i_84;
									for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
										localparam i = _gv_i_84;
										// Trace: src/VX_mem_arb.sv:139:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:140:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 131+:131];
										// Trace: src/VX_mem_arb.sv:141:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_65].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign core_arb.clk = clk;
								assign core_arb.reset = reset;
								genvar _gv_k_1;
								for (_gv_k_1 = 0; _gv_k_1 < NUM_CACHES; _gv_k_1 = _gv_k_1 + 1) begin : g_arb_core_bus_if
									localparam k = _gv_k_1;
									// Trace: src/VX_cache_cluster.sv:83:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].req_valid = arb_core_bus_tmp_if[k].req_valid;
									// Trace: src/VX_cache_cluster.sv:84:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].req_data = arb_core_bus_tmp_if[k].req_data;
									// Trace: src/VX_cache_cluster.sv:85:5
									assign arb_core_bus_tmp_if[k].req_ready = arb_core_bus_if[(k * NUM_REQS) + i].req_ready;
									// Trace: src/VX_cache_cluster.sv:86:5
									assign arb_core_bus_tmp_if[k].rsp_valid = arb_core_bus_if[(k * NUM_REQS) + i].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:87:5
									assign arb_core_bus_tmp_if[k].rsp_data = arb_core_bus_if[(k * NUM_REQS) + i].rsp_data;
									// Trace: src/VX_cache_cluster.sv:88:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].rsp_ready = arb_core_bus_tmp_if[k].rsp_ready;
								end
							end
							// Trace: src/VX_cache_cluster.sv:91:6
							genvar _gv_i_66;
							for (_gv_i_66 = 0; _gv_i_66 < NUM_CACHES; _gv_i_66 = _gv_i_66 + 1) begin : g_cache_wrap
								localparam i = _gv_i_66;
								// Trace: src/VX_cache_cluster.sv:92:9
								// expanded module instance: cache_wrap
								localparam _bbase_665FE_core_bus_if = i * NUM_REQS;
								localparam _bbase_665FE_mem_bus_if = i * MEM_PORTS;
								localparam _param_665FE_INSTANCE_ID = "";
								localparam _param_665FE_CACHE_SIZE = CACHE_SIZE;
								localparam _param_665FE_LINE_SIZE = LINE_SIZE;
								localparam _param_665FE_NUM_BANKS = NUM_BANKS;
								localparam _param_665FE_NUM_WAYS = NUM_WAYS;
								localparam _param_665FE_WORD_SIZE = WORD_SIZE;
								localparam _param_665FE_NUM_REQS = NUM_REQS;
								localparam _param_665FE_MEM_PORTS = MEM_PORTS;
								localparam _param_665FE_WRITE_ENABLE = WRITE_ENABLE;
								localparam _param_665FE_WRITEBACK = WRITEBACK;
								localparam _param_665FE_DIRTY_BYTES = DIRTY_BYTES;
								localparam _param_665FE_REPL_POLICY = REPL_POLICY;
								localparam _param_665FE_CRSQ_SIZE = CRSQ_SIZE;
								localparam _param_665FE_MSHR_SIZE = MSHR_SIZE;
								localparam _param_665FE_MRSQ_SIZE = MRSQ_SIZE;
								localparam _param_665FE_MREQ_SIZE = MREQ_SIZE;
								localparam _param_665FE_UUID_WIDTH = UUID_WIDTH;
								localparam _param_665FE_TAG_WIDTH = ARB_TAG_WIDTH;
								localparam _param_665FE_FLAGS_WIDTH = FLAGS_WIDTH;
								localparam _param_665FE_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_665FE_CORE_OUT_BUF = CORE_OUT_BUF;
								localparam _param_665FE_MEM_OUT_BUF = MEM_OUT_BUF;
								localparam _param_665FE_NC_ENABLE = NC_ENABLE;
								localparam _param_665FE_PASSTHRU = PASSTHRU;
								if (1) begin : cache_wrap
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_cache_wrap.sv:2:16
									localparam INSTANCE_ID = _param_665FE_INSTANCE_ID;
									// Trace: src/VX_cache_wrap.sv:3:15
									localparam TAG_SEL_IDX = _param_665FE_TAG_SEL_IDX;
									// Trace: src/VX_cache_wrap.sv:4:15
									localparam NUM_REQS = _param_665FE_NUM_REQS;
									// Trace: src/VX_cache_wrap.sv:5:15
									localparam MEM_PORTS = _param_665FE_MEM_PORTS;
									// Trace: src/VX_cache_wrap.sv:6:15
									localparam CACHE_SIZE = _param_665FE_CACHE_SIZE;
									// Trace: src/VX_cache_wrap.sv:7:15
									localparam LINE_SIZE = _param_665FE_LINE_SIZE;
									// Trace: src/VX_cache_wrap.sv:8:15
									localparam NUM_BANKS = _param_665FE_NUM_BANKS;
									// Trace: src/VX_cache_wrap.sv:9:15
									localparam NUM_WAYS = _param_665FE_NUM_WAYS;
									// Trace: src/VX_cache_wrap.sv:10:15
									localparam WORD_SIZE = _param_665FE_WORD_SIZE;
									// Trace: src/VX_cache_wrap.sv:11:15
									localparam CRSQ_SIZE = _param_665FE_CRSQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:12:15
									localparam MSHR_SIZE = _param_665FE_MSHR_SIZE;
									// Trace: src/VX_cache_wrap.sv:13:15
									localparam MRSQ_SIZE = _param_665FE_MRSQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:14:15
									localparam MREQ_SIZE = _param_665FE_MREQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:15:15
									localparam WRITE_ENABLE = _param_665FE_WRITE_ENABLE;
									// Trace: src/VX_cache_wrap.sv:16:15
									localparam WRITEBACK = _param_665FE_WRITEBACK;
									// Trace: src/VX_cache_wrap.sv:17:15
									localparam DIRTY_BYTES = _param_665FE_DIRTY_BYTES;
									// Trace: src/VX_cache_wrap.sv:18:15
									localparam REPL_POLICY = _param_665FE_REPL_POLICY;
									// Trace: src/VX_cache_wrap.sv:19:15
									localparam UUID_WIDTH = _param_665FE_UUID_WIDTH;
									// Trace: src/VX_cache_wrap.sv:20:15
									localparam TAG_WIDTH = _param_665FE_TAG_WIDTH;
									// Trace: src/VX_cache_wrap.sv:21:15
									localparam FLAGS_WIDTH = _param_665FE_FLAGS_WIDTH;
									// Trace: src/VX_cache_wrap.sv:22:15
									localparam NC_ENABLE = _param_665FE_NC_ENABLE;
									// Trace: src/VX_cache_wrap.sv:23:15
									localparam PASSTHRU = _param_665FE_PASSTHRU;
									// Trace: src/VX_cache_wrap.sv:24:15
									localparam CORE_OUT_BUF = _param_665FE_CORE_OUT_BUF;
									// Trace: src/VX_cache_wrap.sv:25:15
									localparam MEM_OUT_BUF = _param_665FE_MEM_OUT_BUF;
									// Trace: src/VX_cache_wrap.sv:27:5
									wire clk;
									// Trace: src/VX_cache_wrap.sv:28:5
									wire reset;
									// Trace: src/VX_cache_wrap.sv:29:5
									localparam _mbase_core_bus_if = _bbase_665FE_core_bus_if;
									// Trace: src/VX_cache_wrap.sv:30:5
									localparam _mbase_mem_bus_if = _bbase_665FE_mem_bus_if;
									// Trace: src/VX_cache_wrap.sv:32:5
									localparam CACHE_MEM_TAG_WIDTH = 5;
									// Trace: src/VX_cache_wrap.sv:34:5
									localparam BYPASS_TAG_WIDTH = 5;
									// Trace: src/VX_cache_wrap.sv:36:5
									localparam NC_TAG_WIDTH = 6;
									// Trace: src/VX_cache_wrap.sv:37:5
									localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
									// Trace: src/VX_cache_wrap.sv:38:5
									localparam BYPASS_ENABLE = 1'd1;
									// Trace: src/VX_cache_wrap.sv:39:5
									// expanded interface instance: core_bus_cache_if
									localparam _param_24C1C_DATA_SIZE = WORD_SIZE;
									localparam _param_24C1C_TAG_WIDTH = TAG_WIDTH;
									genvar _arr_24C1C;
									for (_arr_24C1C = 0; _arr_24C1C <= 0; _arr_24C1C = _arr_24C1C + 1) begin : core_bus_cache_if
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_24C1C_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_24C1C_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 28;
										// Trace: src/VX_mem_bus_if.sv:7:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_mem_bus_if.sv:9:5
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:21:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire [178:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire [130:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:30:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:31:5
										// Trace: src/VX_mem_bus_if.sv:39:5
									end
									// Trace: src/VX_cache_wrap.sv:43:5
									// expanded interface instance: mem_bus_cache_if
									localparam _param_D895D_DATA_SIZE = LINE_SIZE;
									localparam _param_D895D_TAG_WIDTH = CACHE_MEM_TAG_WIDTH;
									genvar _arr_D895D;
									for (_arr_D895D = 0; _arr_D895D <= 0; _arr_D895D = _arr_D895D + 1) begin : mem_bus_cache_if
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_D895D_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_D895D_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 26;
										// Trace: src/VX_mem_bus_if.sv:7:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_mem_bus_if.sv:9:5
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:21:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire [610:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire [516:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:30:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:31:5
										// Trace: src/VX_mem_bus_if.sv:39:5
									end
									// Trace: src/VX_cache_wrap.sv:47:5
									// expanded interface instance: mem_bus_tmp_if
									localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
									localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
									genvar _arr_4FE36;
									for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 26;
										// Trace: src/VX_mem_bus_if.sv:7:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_mem_bus_if.sv:9:5
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:21:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire [611:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire [517:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:30:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:31:5
										// Trace: src/VX_mem_bus_if.sv:39:5
									end
									// Trace: src/VX_cache_wrap.sv:51:5
									if (BYPASS_ENABLE) begin : g_bypass
										// Trace: src/VX_cache_wrap.sv:52:9
										// expanded module instance: cache_bypass
										localparam _bbase_714AA_core_bus_in_if = i * NUM_REQS;
										localparam _bbase_714AA_core_bus_out_if = 0;
										localparam _bbase_714AA_mem_bus_in_if = 0;
										localparam _bbase_714AA_mem_bus_out_if = 0;
										localparam _param_714AA_NUM_REQS = NUM_REQS;
										localparam _param_714AA_MEM_PORTS = MEM_PORTS;
										localparam _param_714AA_TAG_SEL_IDX = TAG_SEL_IDX;
										localparam _param_714AA_CACHE_ENABLE = !PASSTHRU;
										localparam _param_714AA_WORD_SIZE = WORD_SIZE;
										localparam _param_714AA_LINE_SIZE = LINE_SIZE;
										localparam _param_714AA_CORE_ADDR_WIDTH = 28;
										localparam _param_714AA_CORE_TAG_WIDTH = TAG_WIDTH;
										localparam _param_714AA_MEM_ADDR_WIDTH = 26;
										localparam _param_714AA_MEM_TAG_IN_WIDTH = CACHE_MEM_TAG_WIDTH;
										localparam _param_714AA_UUID_WIDTH = UUID_WIDTH;
										localparam _param_714AA_CORE_OUT_BUF = CORE_OUT_BUF;
										localparam _param_714AA_MEM_OUT_BUF = MEM_OUT_BUF;
										if (1) begin : cache_bypass
											// Trace: src/VX_cache_bypass.sv:2:15
											localparam NUM_REQS = _param_714AA_NUM_REQS;
											// Trace: src/VX_cache_bypass.sv:3:15
											localparam MEM_PORTS = _param_714AA_MEM_PORTS;
											// Trace: src/VX_cache_bypass.sv:4:15
											localparam TAG_SEL_IDX = _param_714AA_TAG_SEL_IDX;
											// Trace: src/VX_cache_bypass.sv:5:15
											localparam CACHE_ENABLE = _param_714AA_CACHE_ENABLE;
											// Trace: src/VX_cache_bypass.sv:6:15
											localparam WORD_SIZE = _param_714AA_WORD_SIZE;
											// Trace: src/VX_cache_bypass.sv:7:15
											localparam LINE_SIZE = _param_714AA_LINE_SIZE;
											// Trace: src/VX_cache_bypass.sv:8:15
											localparam CORE_ADDR_WIDTH = _param_714AA_CORE_ADDR_WIDTH;
											// Trace: src/VX_cache_bypass.sv:9:15
											localparam CORE_TAG_WIDTH = _param_714AA_CORE_TAG_WIDTH;
											// Trace: src/VX_cache_bypass.sv:10:15
											localparam MEM_ADDR_WIDTH = _param_714AA_MEM_ADDR_WIDTH;
											// Trace: src/VX_cache_bypass.sv:11:15
											localparam MEM_TAG_IN_WIDTH = _param_714AA_MEM_TAG_IN_WIDTH;
											// Trace: src/VX_cache_bypass.sv:12:15
											localparam UUID_WIDTH = _param_714AA_UUID_WIDTH;
											// Trace: src/VX_cache_bypass.sv:13:15
											localparam CORE_OUT_BUF = _param_714AA_CORE_OUT_BUF;
											// Trace: src/VX_cache_bypass.sv:14:15
											localparam MEM_OUT_BUF = _param_714AA_MEM_OUT_BUF;
											// Trace: src/VX_cache_bypass.sv:16:5
											wire clk;
											// Trace: src/VX_cache_bypass.sv:17:5
											wire reset;
											// Trace: src/VX_cache_bypass.sv:18:5
											localparam _mbase_core_bus_in_if = _bbase_714AA_core_bus_in_if;
											// Trace: src/VX_cache_bypass.sv:19:5
											localparam _mbase_core_bus_out_if = 0;
											// Trace: src/VX_cache_bypass.sv:20:5
											localparam _mbase_mem_bus_in_if = 0;
											// Trace: src/VX_cache_bypass.sv:21:5
											localparam _mbase_mem_bus_out_if = 0;
											// Trace: src/VX_cache_bypass.sv:23:5
											localparam DIRECT_PASSTHRU = (!CACHE_ENABLE && 1'd0) && 1'd1;
											// Trace: src/VX_cache_bypass.sv:24:5
											localparam CORE_DATA_WIDTH = 128;
											// Trace: src/VX_cache_bypass.sv:25:5
											localparam WORDS_PER_LINE = 4;
											// Trace: src/VX_cache_bypass.sv:26:5
											localparam WSEL_BITS = 2;
											// Trace: src/VX_cache_bypass.sv:27:5
											localparam CORE_TAG_ID_WIDTH = 2;
											// Trace: src/VX_cache_bypass.sv:28:5
											localparam MEM_TAG_ID_WIDTH = 2;
											// Trace: src/VX_cache_bypass.sv:29:5
											localparam MEM_TAG_NC1_WIDTH = 3;
											// Trace: src/VX_cache_bypass.sv:30:5
											localparam MEM_TAG_NC2_WIDTH = 5;
											// Trace: src/VX_cache_bypass.sv:31:5
											localparam MEM_TAG_OUT_WIDTH = (CACHE_ENABLE ? MEM_TAG_NC2_WIDTH : MEM_TAG_NC2_WIDTH);
											// Trace: src/VX_cache_bypass.sv:32:5
											// expanded interface instance: core_bus_nc_switch_if
											localparam _param_95306_DATA_SIZE = WORD_SIZE;
											localparam _param_95306_TAG_WIDTH = CORE_TAG_WIDTH;
											genvar _arr_95306;
											for (_arr_95306 = 0; _arr_95306 <= (((CACHE_ENABLE ? 2 : 1) * NUM_REQS) - 1); _arr_95306 = _arr_95306 + 1) begin : core_bus_nc_switch_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_95306_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_95306_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [178:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [130:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:36:5
											wire [0:0] core_req_nc_sel;
											// Trace: src/VX_cache_bypass.sv:37:5
											genvar _gv_i_179;
											for (_gv_i_179 = 0; _gv_i_179 < NUM_REQS; _gv_i_179 = _gv_i_179 + 1) begin : g_core_req_is_nc
												localparam i = _gv_i_179;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:39:13
													assign core_req_nc_sel[i] = ~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_in_if].req_data[4];
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:41:13
													assign core_req_nc_sel[i] = 1'b0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:44:5
											// expanded module instance: core_bus_nc_switch
											localparam _bbase_69FDB_bus_in_if = i * NUM_REQS;
											localparam _bbase_69FDB_bus_out_if = 0;
											localparam _param_69FDB_NUM_INPUTS = NUM_REQS;
											localparam _param_69FDB_NUM_OUTPUTS = (CACHE_ENABLE ? 2 : 1) * NUM_REQS;
											localparam _param_69FDB_DATA_SIZE = WORD_SIZE;
											localparam _param_69FDB_TAG_WIDTH = CORE_TAG_WIDTH;
											localparam _param_69FDB_ARBITER = "R";
											localparam _param_69FDB_REQ_OUT_BUF = 0;
											localparam _param_69FDB_RSP_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
											if (1) begin : core_bus_nc_switch
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_switch.sv:2:15
												localparam NUM_INPUTS = _param_69FDB_NUM_INPUTS;
												// Trace: src/VX_mem_switch.sv:3:15
												localparam NUM_OUTPUTS = _param_69FDB_NUM_OUTPUTS;
												// Trace: src/VX_mem_switch.sv:4:15
												localparam DATA_SIZE = _param_69FDB_DATA_SIZE;
												// Trace: src/VX_mem_switch.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_switch.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_switch.sv:7:15
												localparam TAG_WIDTH = _param_69FDB_TAG_WIDTH;
												// Trace: src/VX_mem_switch.sv:8:15
												localparam REQ_OUT_BUF = _param_69FDB_REQ_OUT_BUF;
												// Trace: src/VX_mem_switch.sv:9:15
												localparam RSP_OUT_BUF = _param_69FDB_RSP_OUT_BUF;
												// Trace: src/VX_mem_switch.sv:10:16
												localparam ARBITER = _param_69FDB_ARBITER;
												// Trace: src/VX_mem_switch.sv:11:15
												localparam NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
												// Trace: src/VX_mem_switch.sv:12:15
												localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
												// Trace: src/VX_mem_switch.sv:13:15
												localparam LOG_NUM_REQS = $clog2(NUM_REQS);
												// Trace: src/VX_mem_switch.sv:15:5
												wire clk;
												// Trace: src/VX_mem_switch.sv:16:5
												wire reset;
												// Trace: src/VX_mem_switch.sv:17:5
												wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] bus_sel;
												// Trace: src/VX_mem_switch.sv:18:5
												localparam _mbase_bus_in_if = _bbase_69FDB_bus_in_if;
												// Trace: src/VX_mem_switch.sv:19:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_switch.sv:21:5
												localparam DATA_WIDTH = 128;
												// Trace: src/VX_mem_switch.sv:22:5
												localparam REQ_DATAW = 179;
												// Trace: src/VX_mem_switch.sv:23:5
												localparam RSP_DATAW = 131;
												// Trace: src/VX_mem_switch.sv:24:5
												wire [0:0] req_valid_in;
												// Trace: src/VX_mem_switch.sv:25:5
												wire [178:0] req_data_in;
												// Trace: src/VX_mem_switch.sv:26:5
												wire [0:0] req_ready_in;
												// Trace: src/VX_mem_switch.sv:27:5
												wire [NUM_OUTPUTS - 1:0] req_valid_out;
												// Trace: src/VX_mem_switch.sv:28:5
												wire [(NUM_OUTPUTS * 179) - 1:0] req_data_out;
												// Trace: src/VX_mem_switch.sv:29:5
												wire [NUM_OUTPUTS - 1:0] req_ready_out;
												// Trace: src/VX_mem_switch.sv:30:5
												genvar _gv_i_154;
												for (_gv_i_154 = 0; _gv_i_154 < NUM_INPUTS; _gv_i_154 = _gv_i_154 + 1) begin : g_req_data_in
													localparam i = _gv_i_154;
													// Trace: src/VX_mem_switch.sv:31:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_switch.sv:32:9
													assign req_data_in[i * 179+:179] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_switch.sv:33:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_switch.sv:35:5
												VX_stream_switch #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.OUT_BUF(REQ_OUT_BUF)
												) req_switch(
													.clk(clk),
													.reset(reset),
													.sel_in(bus_sel),
													.valid_in(req_valid_in),
													.data_in(req_data_in),
													.ready_in(req_ready_in),
													.valid_out(req_valid_out),
													.data_out(req_data_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_switch.sv:51:5
												genvar _gv_i_155;
												for (_gv_i_155 = 0; _gv_i_155 < NUM_OUTPUTS; _gv_i_155 = _gv_i_155 + 1) begin : g_req_data_out
													localparam i = _gv_i_155;
													// Trace: src/VX_mem_switch.sv:52:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_switch.sv:53:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_data = req_data_out[i * 179+:179];
													// Trace: src/VX_mem_switch.sv:54:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_ready;
												end
												// Trace: src/VX_mem_switch.sv:56:5
												wire [NUM_OUTPUTS - 1:0] rsp_valid_in;
												// Trace: src/VX_mem_switch.sv:57:5
												wire [(NUM_OUTPUTS * 131) - 1:0] rsp_data_in;
												// Trace: src/VX_mem_switch.sv:58:5
												wire [NUM_OUTPUTS - 1:0] rsp_ready_in;
												// Trace: src/VX_mem_switch.sv:59:5
												wire [0:0] rsp_valid_out;
												// Trace: src/VX_mem_switch.sv:60:5
												wire [130:0] rsp_data_out;
												// Trace: src/VX_mem_switch.sv:61:5
												wire [0:0] rsp_ready_out;
												// Trace: src/VX_mem_switch.sv:62:5
												genvar _gv_i_156;
												for (_gv_i_156 = 0; _gv_i_156 < NUM_OUTPUTS; _gv_i_156 = _gv_i_156 + 1) begin : g_rsp_data_in
													localparam i = _gv_i_156;
													// Trace: src/VX_mem_switch.sv:63:9
													assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_valid;
													// Trace: src/VX_mem_switch.sv:64:9
													assign rsp_data_in[i * 131+:131] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_data;
													// Trace: src/VX_mem_switch.sv:65:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
												end
												// Trace: src/VX_mem_switch.sv:67:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_OUTPUTS),
													.NUM_OUTPUTS(NUM_INPUTS),
													.DATAW(RSP_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(RSP_OUT_BUF)
												) rsp_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(rsp_valid_in),
													.data_in(rsp_data_in),
													.ready_in(rsp_ready_in),
													.valid_out(rsp_valid_out),
													.data_out(rsp_data_out),
													.ready_out(rsp_ready_out),
													.sel_out()
												);
												// Trace: src/VX_mem_switch.sv:84:5
												genvar _gv_i_157;
												for (_gv_i_157 = 0; _gv_i_157 < NUM_INPUTS; _gv_i_157 = _gv_i_157 + 1) begin : g_rsp_data_out
													localparam i = _gv_i_157;
													// Trace: src/VX_mem_switch.sv:85:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_switch.sv:86:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 131+:131];
													// Trace: src/VX_mem_switch.sv:87:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign core_bus_nc_switch.clk = clk;
											assign core_bus_nc_switch.reset = reset;
											assign core_bus_nc_switch.bus_sel = core_req_nc_sel;
											// Trace: src/VX_cache_bypass.sv:59:5
											// expanded interface instance: core_bus_in_nc_if
											localparam _param_C0263_DATA_SIZE = WORD_SIZE;
											localparam _param_C0263_TAG_WIDTH = CORE_TAG_WIDTH;
											genvar _arr_C0263;
											for (_arr_C0263 = 0; _arr_C0263 <= 0; _arr_C0263 = _arr_C0263 + 1) begin : core_bus_in_nc_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_C0263_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_C0263_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [178:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [130:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:63:5
											genvar _gv_i_180;
											for (_gv_i_180 = 0; _gv_i_180 < NUM_REQS; _gv_i_180 = _gv_i_180 + 1) begin : g_core_bus_nc_switch_if
												localparam i = _gv_i_180;
												// Trace: src/VX_cache_bypass.sv:64:9
												assign core_bus_in_nc_if[i].req_valid = core_bus_nc_switch_if[0 + i].req_valid;
												// Trace: src/VX_cache_bypass.sv:65:9
												assign core_bus_in_nc_if[i].req_data = core_bus_nc_switch_if[0 + i].req_data;
												// Trace: src/VX_cache_bypass.sv:66:9
												assign core_bus_nc_switch_if[0 + i].req_ready = core_bus_in_nc_if[i].req_ready;
												// Trace: src/VX_cache_bypass.sv:67:9
												assign core_bus_nc_switch_if[0 + i].rsp_valid = core_bus_in_nc_if[i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:68:9
												assign core_bus_nc_switch_if[0 + i].rsp_data = core_bus_in_nc_if[i].rsp_data;
												// Trace: src/VX_cache_bypass.sv:69:9
												assign core_bus_in_nc_if[i].rsp_ready = core_bus_nc_switch_if[0 + i].rsp_ready;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:71:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = core_bus_nc_switch_if[1 + i].req_valid;
													// Trace: src/VX_cache_bypass.sv:72:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = core_bus_nc_switch_if[1 + i].req_data;
													// Trace: src/VX_cache_bypass.sv:73:13
													assign core_bus_nc_switch_if[1 + i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_ready;
													// Trace: src/VX_cache_bypass.sv:74:13
													assign core_bus_nc_switch_if[1 + i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_valid;
													// Trace: src/VX_cache_bypass.sv:75:13
													assign core_bus_nc_switch_if[1 + i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_data;
													// Trace: src/VX_cache_bypass.sv:76:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = core_bus_nc_switch_if[1 + i].rsp_ready;
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:78:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = 0;
													// Trace: src/VX_cache_bypass.sv:79:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = 1'sb0;
													// Trace: src/VX_cache_bypass.sv:80:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = 0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:83:5
											// expanded interface instance: core_bus_nc_arb_if
											localparam _param_D50AC_DATA_SIZE = WORD_SIZE;
											localparam _param_D50AC_TAG_WIDTH = MEM_TAG_NC1_WIDTH;
											genvar _arr_D50AC;
											for (_arr_D50AC = 0; _arr_D50AC <= 0; _arr_D50AC = _arr_D50AC + 1) begin : core_bus_nc_arb_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_D50AC_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_D50AC_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [178:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [130:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:87:5
											// expanded module instance: core_bus_nc_arb
											localparam _bbase_1376F_bus_in_if = 0;
											localparam _bbase_1376F_bus_out_if = 0;
											localparam _param_1376F_NUM_INPUTS = NUM_REQS;
											localparam _param_1376F_NUM_OUTPUTS = MEM_PORTS;
											localparam _param_1376F_DATA_SIZE = WORD_SIZE;
											localparam _param_1376F_TAG_WIDTH = CORE_TAG_WIDTH;
											localparam _param_1376F_TAG_SEL_IDX = TAG_SEL_IDX;
											localparam _param_1376F_ARBITER = (CACHE_ENABLE ? "P" : "R");
											localparam _param_1376F_REQ_OUT_BUF = 0;
											localparam _param_1376F_RSP_OUT_BUF = 0;
											if (1) begin : core_bus_nc_arb
												// Trace: src/VX_mem_arb.sv:2:15
												localparam NUM_INPUTS = _param_1376F_NUM_INPUTS;
												// Trace: src/VX_mem_arb.sv:3:15
												localparam NUM_OUTPUTS = _param_1376F_NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:4:15
												localparam DATA_SIZE = _param_1376F_DATA_SIZE;
												// Trace: src/VX_mem_arb.sv:5:15
												localparam TAG_WIDTH = _param_1376F_TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:6:15
												localparam TAG_SEL_IDX = _param_1376F_TAG_SEL_IDX;
												// Trace: src/VX_mem_arb.sv:7:15
												localparam REQ_OUT_BUF = _param_1376F_REQ_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:8:15
												localparam RSP_OUT_BUF = _param_1376F_RSP_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:9:16
												localparam ARBITER = _param_1376F_ARBITER;
												// Trace: src/VX_mem_arb.sv:10:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:11:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_arb.sv:12:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_arb.sv:14:5
												wire clk;
												// Trace: src/VX_mem_arb.sv:15:5
												wire reset;
												// Trace: src/VX_mem_arb.sv:16:5
												localparam _mbase_bus_in_if = 0;
												// Trace: src/VX_mem_arb.sv:17:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_arb.sv:19:5
												localparam DATA_WIDTH = 128;
												// Trace: src/VX_mem_arb.sv:20:5
												localparam LOG_NUM_REQS = 0;
												// Trace: src/VX_mem_arb.sv:21:5
												localparam REQ_DATAW = 179;
												// Trace: src/VX_mem_arb.sv:22:5
												localparam RSP_DATAW = 131;
												// Trace: src/VX_mem_arb.sv:24:5
												wire [0:0] req_valid_in;
												// Trace: src/VX_mem_arb.sv:25:5
												wire [178:0] req_data_in;
												// Trace: src/VX_mem_arb.sv:26:5
												wire [0:0] req_ready_in;
												// Trace: src/VX_mem_arb.sv:27:5
												wire [0:0] req_valid_out;
												// Trace: src/VX_mem_arb.sv:28:5
												wire [178:0] req_data_out;
												// Trace: src/VX_mem_arb.sv:29:5
												wire [0:0] req_sel_out;
												// Trace: src/VX_mem_arb.sv:30:5
												wire [0:0] req_ready_out;
												// Trace: src/VX_mem_arb.sv:31:5
												genvar _gv_i_80;
												for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
													localparam i = _gv_i_80;
													// Trace: src/VX_mem_arb.sv:32:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_arb.sv:33:9
													assign req_data_in[i * 179+:179] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_arb.sv:34:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_arb.sv:36:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(REQ_OUT_BUF)
												) req_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(req_valid_in),
													.ready_in(req_ready_in),
													.data_in(req_data_in),
													.data_out(req_data_out),
													.sel_out(req_sel_out),
													.valid_out(req_valid_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_arb.sv:53:5
												genvar _gv_i_81;
												for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
													localparam i = _gv_i_81;
													// Trace: src/VX_mem_arb.sv:54:9
													wire [2:0] req_tag_out;
													// Trace: src/VX_mem_arb.sv:55:9
													VX_bits_insert #(
														.N(TAG_WIDTH),
														.S(LOG_NUM_REQS),
														.POS(TAG_SEL_IDX)
													) bits_insert(
														.data_in(req_tag_out),
														.ins_in(req_sel_out[i+:1]),
														.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[2-:3])
													);
													// Trace: src/VX_mem_arb.sv:64:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_arb.sv:65:9
													assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[178], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[177-:28], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[149-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[21-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[5-:3], req_tag_out} = req_data_out[i * 179+:179];
													// Trace: src/VX_mem_arb.sv:73:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_ready;
												end
												// Trace: src/VX_mem_arb.sv:75:5
												wire [0:0] rsp_valid_out;
												// Trace: src/VX_mem_arb.sv:76:5
												wire [130:0] rsp_data_out;
												// Trace: src/VX_mem_arb.sv:77:5
												wire [0:0] rsp_ready_out;
												// Trace: src/VX_mem_arb.sv:78:5
												wire [0:0] rsp_valid_in;
												// Trace: src/VX_mem_arb.sv:79:5
												wire [130:0] rsp_data_in;
												// Trace: src/VX_mem_arb.sv:80:5
												wire [0:0] rsp_ready_in;
												// Trace: src/VX_mem_arb.sv:81:5
												if (1) begin : g_passthru
													genvar _gv_i_83;
													for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_83;
														// Trace: src/VX_mem_arb.sv:116:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:117:13
														assign rsp_data_in[i * 131+:131] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_data;
														// Trace: src/VX_mem_arb.sv:118:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:120:9
													VX_stream_arb #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.ARBITER(ARBITER),
														.OUT_BUF(RSP_OUT_BUF)
													) req_arb(
														.clk(clk),
														.reset(reset),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out),
														.sel_out()
													);
												end
												// Trace: src/VX_mem_arb.sv:138:5
												genvar _gv_i_84;
												for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
													localparam i = _gv_i_84;
													// Trace: src/VX_mem_arb.sv:139:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_arb.sv:140:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 131+:131];
													// Trace: src/VX_mem_arb.sv:141:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign core_bus_nc_arb.clk = clk;
											assign core_bus_nc_arb.reset = reset;
											// Trace: src/VX_cache_bypass.sv:102:5
											// expanded interface instance: mem_bus_out_nc_if
											localparam _param_0061C_DATA_SIZE = LINE_SIZE;
											localparam _param_0061C_TAG_WIDTH = MEM_TAG_NC2_WIDTH;
											genvar _arr_0061C;
											for (_arr_0061C = 0; _arr_0061C <= 0; _arr_0061C = _arr_0061C + 1) begin : mem_bus_out_nc_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_0061C_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_0061C_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [610:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [516:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:106:5
											genvar _gv_i_181;
											for (_gv_i_181 = 0; _gv_i_181 < MEM_PORTS; _gv_i_181 = _gv_i_181 + 1) begin : g_mem_bus_out_nc
												localparam i = _gv_i_181;
												// Trace: src/VX_cache_bypass.sv:107:9
												wire core_req_nc_arb_rw;
												// Trace: src/VX_cache_bypass.sv:108:9
												wire [15:0] core_req_nc_arb_byteen;
												// Trace: src/VX_cache_bypass.sv:109:9
												wire [27:0] core_req_nc_arb_addr;
												// Trace: src/VX_cache_bypass.sv:110:9
												wire [2:0] core_req_nc_arb_flags;
												// Trace: src/VX_cache_bypass.sv:111:9
												wire [127:0] core_req_nc_arb_data;
												// Trace: src/VX_cache_bypass.sv:112:9
												wire [2:0] core_req_nc_arb_tag;
												// Trace: src/VX_cache_bypass.sv:113:9
												assign {core_req_nc_arb_rw, core_req_nc_arb_addr, core_req_nc_arb_data, core_req_nc_arb_byteen, core_req_nc_arb_flags, core_req_nc_arb_tag} = core_bus_nc_arb_if[i].req_data;
												// Trace: src/VX_cache_bypass.sv:121:9
												wire [25:0] core_req_nc_arb_addr_w;
												// Trace: src/VX_cache_bypass.sv:122:9
												reg [63:0] core_req_nc_arb_byteen_w;
												// Trace: src/VX_cache_bypass.sv:123:9
												reg [511:0] core_req_nc_arb_data_w;
												// Trace: src/VX_cache_bypass.sv:124:9
												wire [127:0] core_rsp_nc_arb_data_w;
												// Trace: src/VX_cache_bypass.sv:125:9
												wire [4:0] core_req_nc_arb_tag_w;
												// Trace: src/VX_cache_bypass.sv:126:9
												wire [2:0] core_rsp_nc_arb_tag_w;
												if (1) begin : g_multi_word_line
													// Trace: src/VX_cache_bypass.sv:128:13
													wire [1:0] rsp_wsel;
													// Trace: src/VX_cache_bypass.sv:129:13
													wire [1:0] req_wsel = core_req_nc_arb_addr[1:0];
													// Trace: src/VX_cache_bypass.sv:130:13
													always @(*) begin
														// Trace: src/VX_cache_bypass.sv:131:17
														core_req_nc_arb_byteen_w = 1'sb0;
														// Trace: src/VX_cache_bypass.sv:132:17
														core_req_nc_arb_byteen_w[req_wsel * 16+:16] = core_req_nc_arb_byteen;
														// Trace: src/VX_cache_bypass.sv:133:17
														core_req_nc_arb_data_w = 1'sbx;
														// Trace: src/VX_cache_bypass.sv:134:17
														core_req_nc_arb_data_w[req_wsel * 128+:128] = core_req_nc_arb_data;
													end
													// Trace: src/VX_cache_bypass.sv:136:13
													VX_bits_insert #(
														.N(MEM_TAG_NC1_WIDTH),
														.S(WSEL_BITS),
														.POS(TAG_SEL_IDX)
													) wsel_insert(
														.data_in(core_req_nc_arb_tag),
														.ins_in(req_wsel),
														.data_out(core_req_nc_arb_tag_w)
													);
													// Trace: src/VX_cache_bypass.sv:145:13
													VX_bits_remove #(
														.N(MEM_TAG_NC2_WIDTH),
														.S(WSEL_BITS),
														.POS(TAG_SEL_IDX)
													) wsel_remove(
														.data_in(mem_bus_out_nc_if[i].rsp_data[4-:5]),
														.sel_out(rsp_wsel),
														.data_out(core_rsp_nc_arb_tag_w)
													);
													// Trace: src/VX_cache_bypass.sv:154:13
													assign core_req_nc_arb_addr_w = core_req_nc_arb_addr[WSEL_BITS+:MEM_ADDR_WIDTH];
													// Trace: src/VX_cache_bypass.sv:155:13
													assign core_rsp_nc_arb_data_w = mem_bus_out_nc_if[i].rsp_data[5 + (rsp_wsel * CORE_DATA_WIDTH)+:CORE_DATA_WIDTH];
												end
												// Trace: src/VX_cache_bypass.sv:164:9
												assign mem_bus_out_nc_if[i].req_valid = core_bus_nc_arb_if[i].req_valid;
												// Trace: src/VX_cache_bypass.sv:165:9
												assign mem_bus_out_nc_if[i].req_data = {core_req_nc_arb_rw, core_req_nc_arb_addr_w, core_req_nc_arb_data_w, core_req_nc_arb_byteen_w, core_req_nc_arb_flags, core_req_nc_arb_tag_w};
												// Trace: src/VX_cache_bypass.sv:173:9
												assign core_bus_nc_arb_if[i].req_ready = mem_bus_out_nc_if[i].req_ready;
												// Trace: src/VX_cache_bypass.sv:174:9
												assign core_bus_nc_arb_if[i].rsp_valid = mem_bus_out_nc_if[i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:175:9
												assign core_bus_nc_arb_if[i].rsp_data = {core_rsp_nc_arb_data_w, core_rsp_nc_arb_tag_w};
												// Trace: src/VX_cache_bypass.sv:179:9
												assign mem_bus_out_nc_if[i].rsp_ready = core_bus_nc_arb_if[i].rsp_ready;
											end
											// Trace: src/VX_cache_bypass.sv:181:5
											// expanded interface instance: mem_bus_out_src_if
											localparam _param_913F6_DATA_SIZE = LINE_SIZE;
											localparam _param_913F6_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
											genvar _arr_913F6;
											for (_arr_913F6 = 0; _arr_913F6 <= (((CACHE_ENABLE ? 2 : 1) * MEM_PORTS) - 1); _arr_913F6 = _arr_913F6 + 1) begin : mem_bus_out_src_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_913F6_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_913F6_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [610:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [516:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache_bypass.sv:185:5
											genvar _gv_i_182;
											for (_gv_i_182 = 0; _gv_i_182 < MEM_PORTS; _gv_i_182 = _gv_i_182 + 1) begin : g_mem_bus_out_src
												localparam i = _gv_i_182;
												// Trace: src/VX_cache_bypass.sv:186:5
												assign mem_bus_out_src_if[0 + i].req_valid = mem_bus_out_nc_if[i].req_valid;
												// Trace: src/VX_cache_bypass.sv:187:5
												assign mem_bus_out_src_if[0 + i].req_data[610] = mem_bus_out_nc_if[i].req_data[610];
												// Trace: src/VX_cache_bypass.sv:188:5
												assign mem_bus_out_src_if[0 + i].req_data[609-:26] = mem_bus_out_nc_if[i].req_data[609-:26];
												// Trace: src/VX_cache_bypass.sv:189:5
												assign mem_bus_out_src_if[0 + i].req_data[583-:512] = mem_bus_out_nc_if[i].req_data[583-:512];
												// Trace: src/VX_cache_bypass.sv:190:5
												assign mem_bus_out_src_if[0 + i].req_data[71-:64] = mem_bus_out_nc_if[i].req_data[71-:64];
												// Trace: src/VX_cache_bypass.sv:191:5
												assign mem_bus_out_src_if[0 + i].req_data[7-:3] = mem_bus_out_nc_if[i].req_data[7-:3];
												if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk1
													if (1) begin : genblk1
														if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
															// Trace: src/VX_cache_bypass.sv:196:17
															assign mem_bus_out_src_if[0 + i].req_data[4-:5] = {mem_bus_out_nc_if[i].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_NC2_WIDTH {1'b0}}, mem_bus_out_nc_if[i].req_data[3-:4]};
														end
														else begin : genblk1
															// Trace: src/VX_cache_bypass.sv:198:17
															assign mem_bus_out_src_if[0 + i].req_data[4-:5] = {mem_bus_out_nc_if[i].req_data[4-:1], mem_bus_out_nc_if[i].req_data[(MEM_TAG_OUT_WIDTH - UUID_WIDTH) - 1:0]};
														end
													end
												end
												else begin : genblk1
													// Trace: src/VX_cache_bypass.sv:208:9
													assign mem_bus_out_src_if[0 + i].req_data[4-:5] = mem_bus_out_nc_if[i].req_data[4-:5];
												end
												// Trace: src/VX_cache_bypass.sv:211:5
												assign mem_bus_out_nc_if[i].req_ready = mem_bus_out_src_if[0 + i].req_ready;
												// Trace: src/VX_cache_bypass.sv:212:5
												assign mem_bus_out_nc_if[i].rsp_valid = mem_bus_out_src_if[0 + i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:213:5
												assign mem_bus_out_nc_if[i].rsp_data[516-:512] = mem_bus_out_src_if[0 + i].rsp_data[516-:512];
												if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk2
													if (1) begin : genblk1
														if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
															// Trace: src/VX_cache_bypass.sv:218:17
															assign mem_bus_out_nc_if[i].rsp_data[4-:5] = {mem_bus_out_src_if[0 + i].rsp_data[4-:1], mem_bus_out_src_if[0 + i].rsp_data[3:0]};
														end
														else begin : genblk1
															// Trace: src/VX_cache_bypass.sv:220:17
															assign mem_bus_out_nc_if[i].rsp_data[4-:5] = {mem_bus_out_src_if[0 + i].rsp_data[4-:1], {MEM_TAG_NC2_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[0 + i].rsp_data[3-:4]};
														end
													end
												end
												else begin : genblk2
													// Trace: src/VX_cache_bypass.sv:230:9
													assign mem_bus_out_nc_if[i].rsp_data[4-:5] = mem_bus_out_src_if[0 + i].rsp_data[4-:5];
												end
												// Trace: src/VX_cache_bypass.sv:233:5
												assign mem_bus_out_src_if[0 + i].rsp_ready = mem_bus_out_nc_if[i].rsp_ready;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:235:5
													assign mem_bus_out_src_if[1 + i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_valid;
													// Trace: src/VX_cache_bypass.sv:236:5
													assign mem_bus_out_src_if[1 + i].req_data[610] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[610];
													// Trace: src/VX_cache_bypass.sv:237:5
													assign mem_bus_out_src_if[1 + i].req_data[609-:26] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[609-:26];
													// Trace: src/VX_cache_bypass.sv:238:5
													assign mem_bus_out_src_if[1 + i].req_data[583-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[583-:512];
													// Trace: src/VX_cache_bypass.sv:239:5
													assign mem_bus_out_src_if[1 + i].req_data[71-:64] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[71-:64];
													// Trace: src/VX_cache_bypass.sv:240:5
													assign mem_bus_out_src_if[1 + i].req_data[7-:3] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[7-:3];
													if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk1
														if (1) begin : genblk1
															if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
																// Trace: src/VX_cache_bypass.sv:245:17
																assign mem_bus_out_src_if[1 + i].req_data[4-:5] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_IN_WIDTH {1'b0}}, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[3-:4]};
															end
															else begin : genblk1
																// Trace: src/VX_cache_bypass.sv:247:17
																assign mem_bus_out_src_if[1 + i].req_data[4-:5] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[(MEM_TAG_OUT_WIDTH - UUID_WIDTH) - 1:0]};
															end
														end
													end
													else begin : genblk1
														// Trace: src/VX_cache_bypass.sv:257:9
														assign mem_bus_out_src_if[1 + i].req_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:5];
													end
													// Trace: src/VX_cache_bypass.sv:260:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = mem_bus_out_src_if[1 + i].req_ready;
													// Trace: src/VX_cache_bypass.sv:261:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = mem_bus_out_src_if[1 + i].rsp_valid;
													// Trace: src/VX_cache_bypass.sv:262:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[516-:512] = mem_bus_out_src_if[1 + i].rsp_data[516-:512];
													if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk2
														if (1) begin : genblk1
															if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
																// Trace: src/VX_cache_bypass.sv:267:17
																assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[4-:1], mem_bus_out_src_if[1 + i].rsp_data[3:0]};
															end
															else begin : genblk1
																// Trace: src/VX_cache_bypass.sv:269:17
																assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[4-:1], {MEM_TAG_IN_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[1 + i].rsp_data[3-:4]};
															end
														end
													end
													else begin : genblk2
														// Trace: src/VX_cache_bypass.sv:279:9
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = mem_bus_out_src_if[1 + i].rsp_data[4-:5];
													end
													// Trace: src/VX_cache_bypass.sv:282:5
													assign mem_bus_out_src_if[1 + i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_ready;
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:284:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = 0;
													// Trace: src/VX_cache_bypass.sv:285:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = 0;
													// Trace: src/VX_cache_bypass.sv:286:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data = 1'sb0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:289:5
											// expanded module instance: mem_bus_out_arb
											localparam _bbase_B06D0_bus_in_if = 0;
											localparam _bbase_B06D0_bus_out_if = 0;
											localparam _param_B06D0_NUM_INPUTS = (CACHE_ENABLE ? 2 : 1) * MEM_PORTS;
											localparam _param_B06D0_NUM_OUTPUTS = MEM_PORTS;
											localparam _param_B06D0_DATA_SIZE = LINE_SIZE;
											localparam _param_B06D0_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
											localparam _param_B06D0_ARBITER = "R";
											localparam _param_B06D0_REQ_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
											localparam _param_B06D0_RSP_OUT_BUF = 0;
											if (1) begin : mem_bus_out_arb
												// Trace: src/VX_mem_arb.sv:2:15
												localparam NUM_INPUTS = _param_B06D0_NUM_INPUTS;
												// Trace: src/VX_mem_arb.sv:3:15
												localparam NUM_OUTPUTS = _param_B06D0_NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:4:15
												localparam DATA_SIZE = _param_B06D0_DATA_SIZE;
												// Trace: src/VX_mem_arb.sv:5:15
												localparam TAG_WIDTH = _param_B06D0_TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:6:15
												localparam TAG_SEL_IDX = 0;
												// Trace: src/VX_mem_arb.sv:7:15
												localparam REQ_OUT_BUF = _param_B06D0_REQ_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:8:15
												localparam RSP_OUT_BUF = _param_B06D0_RSP_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:9:16
												localparam ARBITER = _param_B06D0_ARBITER;
												// Trace: src/VX_mem_arb.sv:10:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:11:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_arb.sv:12:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_arb.sv:14:5
												wire clk;
												// Trace: src/VX_mem_arb.sv:15:5
												wire reset;
												// Trace: src/VX_mem_arb.sv:16:5
												localparam _mbase_bus_in_if = 0;
												// Trace: src/VX_mem_arb.sv:17:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_arb.sv:19:5
												localparam DATA_WIDTH = 512;
												// Trace: src/VX_mem_arb.sv:20:5
												localparam LOG_NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? $clog2((NUM_INPUTS + 0) / 1) : 0);
												// Trace: src/VX_mem_arb.sv:21:5
												localparam REQ_DATAW = 606 + TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:22:5
												localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:24:5
												wire [NUM_INPUTS - 1:0] req_valid_in;
												// Trace: src/VX_mem_arb.sv:25:5
												wire [(NUM_INPUTS * REQ_DATAW) - 1:0] req_data_in;
												// Trace: src/VX_mem_arb.sv:26:5
												wire [NUM_INPUTS - 1:0] req_ready_in;
												// Trace: src/VX_mem_arb.sv:27:5
												wire [0:0] req_valid_out;
												// Trace: src/VX_mem_arb.sv:28:5
												wire [REQ_DATAW - 1:0] req_data_out;
												// Trace: src/VX_mem_arb.sv:29:5
												wire [(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1) - 1:0] req_sel_out;
												// Trace: src/VX_mem_arb.sv:30:5
												wire [0:0] req_ready_out;
												// Trace: src/VX_mem_arb.sv:31:5
												genvar _gv_i_80;
												for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
													localparam i = _gv_i_80;
													// Trace: src/VX_mem_arb.sv:32:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_arb.sv:33:9
													assign req_data_in[i * 611+:611] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_arb.sv:34:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_arb.sv:36:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(REQ_OUT_BUF)
												) req_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(req_valid_in),
													.ready_in(req_ready_in),
													.data_in(req_data_in),
													.data_out(req_data_out),
													.sel_out(req_sel_out),
													.valid_out(req_valid_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_arb.sv:53:5
												genvar _gv_i_81;
												for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
													localparam i = _gv_i_81;
													// Trace: src/VX_mem_arb.sv:54:9
													wire [TAG_WIDTH - 1:0] req_tag_out;
													// Trace: src/VX_mem_arb.sv:55:9
													VX_bits_insert #(
														.N(TAG_WIDTH),
														.S(LOG_NUM_REQS),
														.POS(TAG_SEL_IDX)
													) bits_insert(
														.data_in(req_tag_out),
														.ins_in(req_sel_out[i * 1+:1]),
														.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[5-:6])
													);
													// Trace: src/VX_mem_arb.sv:64:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_arb.sv:65:9
													assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[611], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[610-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[584-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[72-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[8-:3], req_tag_out} = req_data_out[i * 611+:611];
													// Trace: src/VX_mem_arb.sv:73:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
												end
												// Trace: src/VX_mem_arb.sv:75:5
												wire [NUM_INPUTS - 1:0] rsp_valid_out;
												// Trace: src/VX_mem_arb.sv:76:5
												wire [(NUM_INPUTS * RSP_DATAW) - 1:0] rsp_data_out;
												// Trace: src/VX_mem_arb.sv:77:5
												wire [NUM_INPUTS - 1:0] rsp_ready_out;
												// Trace: src/VX_mem_arb.sv:78:5
												wire [0:0] rsp_valid_in;
												// Trace: src/VX_mem_arb.sv:79:5
												wire [RSP_DATAW - 1:0] rsp_data_in;
												// Trace: src/VX_mem_arb.sv:80:5
												wire [0:0] rsp_ready_in;
												// Trace: src/VX_mem_arb.sv:81:5
												if (NUM_INPUTS > NUM_OUTPUTS) begin : g_rsp_enabled
													// Trace: src/VX_mem_arb.sv:82:9
													wire [LOG_NUM_REQS - 1:0] rsp_sel_in;
													genvar _gv_i_82;
													for (_gv_i_82 = 0; _gv_i_82 < NUM_OUTPUTS; _gv_i_82 = _gv_i_82 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_82;
														// Trace: src/VX_mem_arb.sv:84:13
														wire [TAG_WIDTH - 1:0] rsp_tag_out;
														// Trace: src/VX_mem_arb.sv:85:13
														VX_bits_remove #(
															.N(TAG_WIDTH + LOG_NUM_REQS),
															.S(LOG_NUM_REQS),
															.POS(TAG_SEL_IDX)
														) bits_remove(
															.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[5-:6]),
															.sel_out(rsp_sel_in[i * 1+:1]),
															.data_out(rsp_tag_out)
														);
														// Trace: src/VX_mem_arb.sv:94:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:95:13
														assign rsp_data_in[i * 517+:517] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[517-:512], rsp_tag_out};
														// Trace: src/VX_mem_arb.sv:96:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:98:9
													VX_stream_switch #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.OUT_BUF(RSP_OUT_BUF)
													) rsp_switch(
														.clk(clk),
														.reset(reset),
														.sel_in(rsp_sel_in),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out)
													);
												end
												else begin : g_passthru
													genvar _gv_i_83;
													for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_83;
														// Trace: src/VX_mem_arb.sv:116:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:117:13
														assign rsp_data_in[i * 517+:517] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
														// Trace: src/VX_mem_arb.sv:118:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:120:9
													VX_stream_arb #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.ARBITER(ARBITER),
														.OUT_BUF(RSP_OUT_BUF)
													) req_arb(
														.clk(clk),
														.reset(reset),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out),
														.sel_out()
													);
												end
												// Trace: src/VX_mem_arb.sv:138:5
												genvar _gv_i_84;
												for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
													localparam i = _gv_i_84;
													// Trace: src/VX_mem_arb.sv:139:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_arb.sv:140:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 517+:517];
													// Trace: src/VX_mem_arb.sv:141:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign mem_bus_out_arb.clk = clk;
											assign mem_bus_out_arb.reset = reset;
										end
										assign cache_bypass.clk = clk;
										assign cache_bypass.reset = reset;
									end
									else begin : g_no_bypass
										genvar _gv_i_167;
										for (_gv_i_167 = 0; _gv_i_167 < NUM_REQS; _gv_i_167 = _gv_i_167 + 1) begin : g_core_bus_cache_if
											localparam i = _gv_i_167;
											// Trace: src/VX_cache_wrap.sv:76:5
											assign core_bus_cache_if[i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].req_valid;
											// Trace: src/VX_cache_wrap.sv:77:5
											assign core_bus_cache_if[i].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].req_data;
											// Trace: src/VX_cache_wrap.sv:78:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].req_ready = core_bus_cache_if[i].req_ready;
											// Trace: src/VX_cache_wrap.sv:79:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_valid = core_bus_cache_if[i].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:80:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_data = core_bus_cache_if[i].rsp_data;
											// Trace: src/VX_cache_wrap.sv:81:5
											assign core_bus_cache_if[i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_ready;
										end
										genvar _gv_i_168;
										for (_gv_i_168 = 0; _gv_i_168 < MEM_PORTS; _gv_i_168 = _gv_i_168 + 1) begin : g_mem_bus_tmp_if
											localparam i = _gv_i_168;
											// Trace: src/VX_cache_wrap.sv:84:5
											assign mem_bus_tmp_if[i].req_valid = mem_bus_cache_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:85:5
											assign mem_bus_tmp_if[i].req_data = mem_bus_cache_if[i].req_data;
											// Trace: src/VX_cache_wrap.sv:86:5
											assign mem_bus_cache_if[i].req_ready = mem_bus_tmp_if[i].req_ready;
											// Trace: src/VX_cache_wrap.sv:87:5
											assign mem_bus_cache_if[i].rsp_valid = mem_bus_tmp_if[i].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:88:5
											assign mem_bus_cache_if[i].rsp_data = mem_bus_tmp_if[i].rsp_data;
											// Trace: src/VX_cache_wrap.sv:89:5
											assign mem_bus_tmp_if[i].rsp_ready = mem_bus_cache_if[i].rsp_ready;
										end
									end
									// Trace: src/VX_cache_wrap.sv:92:5
									genvar _gv_i_169;
									for (_gv_i_169 = 0; _gv_i_169 < MEM_PORTS; _gv_i_169 = _gv_i_169 + 1) begin : g_mem_bus_if
										localparam i = _gv_i_169;
										if (WRITE_ENABLE) begin : g_we
											// Trace: src/VX_cache_wrap.sv:94:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:95:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
											// Trace: src/VX_cache_wrap.sv:96:5
											assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
											// Trace: src/VX_cache_wrap.sv:97:5
											assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:98:5
											assign mem_bus_tmp_if[i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
											// Trace: src/VX_cache_wrap.sv:99:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
										end
										else begin : g_ro
											// Trace: src/VX_cache_wrap.sv:101:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:102:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[611] = 0;
											// Trace: src/VX_cache_wrap.sv:103:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[610-:26] = mem_bus_tmp_if[i].req_data[610-:26];
											// Trace: src/VX_cache_wrap.sv:104:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[584-:512] = 1'sb0;
											// Trace: src/VX_cache_wrap.sv:105:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[72-:64] = 1'sb1;
											// Trace: src/VX_cache_wrap.sv:106:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[8-:3] = mem_bus_tmp_if[i].req_data[8-:3];
											// Trace: src/VX_cache_wrap.sv:107:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[5-:6] = mem_bus_tmp_if[i].req_data[5-:6];
											// Trace: src/VX_cache_wrap.sv:108:5
											assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
											// Trace: src/VX_cache_wrap.sv:109:5
											assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:110:5
											assign mem_bus_tmp_if[i].rsp_data[517-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[517-:512];
											// Trace: src/VX_cache_wrap.sv:111:5
											assign mem_bus_tmp_if[i].rsp_data[5-:6] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[5-:6];
											// Trace: src/VX_cache_wrap.sv:112:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
										end
									end
									// Trace: src/VX_cache_wrap.sv:115:5
									if (1) begin : g_cache
										// Trace: src/VX_cache_wrap.sv:116:9
										// expanded module instance: cache
										localparam _bbase_90EE2_core_bus_if = 0;
										localparam _bbase_90EE2_mem_bus_if = 0;
										localparam _param_90EE2_INSTANCE_ID = INSTANCE_ID;
										localparam _param_90EE2_CACHE_SIZE = CACHE_SIZE;
										localparam _param_90EE2_LINE_SIZE = LINE_SIZE;
										localparam _param_90EE2_NUM_BANKS = NUM_BANKS;
										localparam _param_90EE2_NUM_WAYS = NUM_WAYS;
										localparam _param_90EE2_WORD_SIZE = WORD_SIZE;
										localparam _param_90EE2_NUM_REQS = NUM_REQS;
										localparam _param_90EE2_MEM_PORTS = MEM_PORTS;
										localparam _param_90EE2_WRITE_ENABLE = WRITE_ENABLE;
										localparam _param_90EE2_WRITEBACK = WRITEBACK;
										localparam _param_90EE2_DIRTY_BYTES = DIRTY_BYTES;
										localparam _param_90EE2_REPL_POLICY = REPL_POLICY;
										localparam _param_90EE2_CRSQ_SIZE = CRSQ_SIZE;
										localparam _param_90EE2_MSHR_SIZE = MSHR_SIZE;
										localparam _param_90EE2_MRSQ_SIZE = MRSQ_SIZE;
										localparam _param_90EE2_MREQ_SIZE = MREQ_SIZE;
										localparam _param_90EE2_UUID_WIDTH = UUID_WIDTH;
										localparam _param_90EE2_TAG_WIDTH = TAG_WIDTH;
										localparam _param_90EE2_FLAGS_WIDTH = FLAGS_WIDTH;
										localparam _param_90EE2_CORE_OUT_BUF = (BYPASS_ENABLE ? 1 : CORE_OUT_BUF);
										localparam _param_90EE2_MEM_OUT_BUF = (BYPASS_ENABLE ? 1 : MEM_OUT_BUF);
										if (1) begin : cache
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_cache.sv:2:16
											localparam INSTANCE_ID = _param_90EE2_INSTANCE_ID;
											// Trace: src/VX_cache.sv:3:15
											localparam NUM_REQS = _param_90EE2_NUM_REQS;
											// Trace: src/VX_cache.sv:4:15
											localparam MEM_PORTS = _param_90EE2_MEM_PORTS;
											// Trace: src/VX_cache.sv:5:15
											localparam CACHE_SIZE = _param_90EE2_CACHE_SIZE;
											// Trace: src/VX_cache.sv:6:15
											localparam LINE_SIZE = _param_90EE2_LINE_SIZE;
											// Trace: src/VX_cache.sv:7:15
											localparam NUM_BANKS = _param_90EE2_NUM_BANKS;
											// Trace: src/VX_cache.sv:8:15
											localparam NUM_WAYS = _param_90EE2_NUM_WAYS;
											// Trace: src/VX_cache.sv:9:15
											localparam WORD_SIZE = _param_90EE2_WORD_SIZE;
											// Trace: src/VX_cache.sv:10:15
											localparam CRSQ_SIZE = _param_90EE2_CRSQ_SIZE;
											// Trace: src/VX_cache.sv:11:15
											localparam MSHR_SIZE = _param_90EE2_MSHR_SIZE;
											// Trace: src/VX_cache.sv:12:15
											localparam MRSQ_SIZE = _param_90EE2_MRSQ_SIZE;
											// Trace: src/VX_cache.sv:13:15
											localparam MREQ_SIZE = _param_90EE2_MREQ_SIZE;
											// Trace: src/VX_cache.sv:14:15
											localparam WRITE_ENABLE = _param_90EE2_WRITE_ENABLE;
											// Trace: src/VX_cache.sv:15:15
											localparam WRITEBACK = _param_90EE2_WRITEBACK;
											// Trace: src/VX_cache.sv:16:15
											localparam DIRTY_BYTES = _param_90EE2_DIRTY_BYTES;
											// Trace: src/VX_cache.sv:17:15
											localparam REPL_POLICY = _param_90EE2_REPL_POLICY;
											// Trace: src/VX_cache.sv:18:15
											localparam UUID_WIDTH = _param_90EE2_UUID_WIDTH;
											// Trace: src/VX_cache.sv:19:15
											localparam TAG_WIDTH = _param_90EE2_TAG_WIDTH;
											// Trace: src/VX_cache.sv:20:15
											localparam FLAGS_WIDTH = _param_90EE2_FLAGS_WIDTH;
											// Trace: src/VX_cache.sv:21:15
											localparam CORE_OUT_BUF = _param_90EE2_CORE_OUT_BUF;
											// Trace: src/VX_cache.sv:22:15
											localparam MEM_OUT_BUF = _param_90EE2_MEM_OUT_BUF;
											// Trace: src/VX_cache.sv:24:5
											wire clk;
											// Trace: src/VX_cache.sv:25:5
											wire reset;
											// Trace: src/VX_cache.sv:26:5
											localparam _mbase_core_bus_if = 0;
											// Trace: src/VX_cache.sv:27:5
											localparam _mbase_mem_bus_if = 0;
											// Trace: src/VX_cache.sv:29:5
											localparam REQ_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:30:5
											localparam WORD_SEL_WIDTH = 2;
											// Trace: src/VX_cache.sv:31:5
											localparam MSHR_ADDR_WIDTH = 4;
											// Trace: src/VX_cache.sv:32:5
											localparam MEM_TAG_WIDTH = 5;
											// Trace: src/VX_cache.sv:34:5
											localparam WORDS_PER_LINE = 4;
											// Trace: src/VX_cache.sv:35:5
											localparam WORD_WIDTH = 128;
											// Trace: src/VX_cache.sv:36:5
											localparam WORD_SEL_BITS = 2;
											// Trace: src/VX_cache.sv:37:5
											localparam BANK_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:38:5
											localparam BANK_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:39:5
											localparam LINE_ADDR_WIDTH = 26;
											// Trace: src/VX_cache.sv:40:5
											localparam CORE_REQ_DATAW = 179;
											// Trace: src/VX_cache.sv:41:5
											localparam CORE_RSP_DATAW = 131;
											// Trace: src/VX_cache.sv:42:5
											localparam BANK_MEM_TAG_WIDTH = 5;
											// Trace: src/VX_cache.sv:43:5
											localparam MEM_REQ_DATAW = 611;
											// Trace: src/VX_cache.sv:44:5
											localparam MEM_RSP_DATAW = 517;
											// Trace: src/VX_cache.sv:45:5
											localparam MEM_PORTS_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:46:5
											localparam MEM_PORTS_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:47:5
											localparam MEM_ARB_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:48:5
											localparam MEM_ARB_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:49:5
											localparam CORE_RSP_REG_DISABLE = 1'd0;
											// Trace: src/VX_cache.sv:50:5
											localparam MEM_REQ_REG_DISABLE = 1'd0;
											// Trace: src/VX_cache.sv:51:5
											localparam REQ_XBAR_BUF = 0;
											// Trace: src/VX_cache.sv:52:5
											// expanded interface instance: core_bus2_if
											localparam _param_9260A_DATA_SIZE = WORD_SIZE;
											localparam _param_9260A_TAG_WIDTH = TAG_WIDTH;
											genvar _arr_9260A;
											for (_arr_9260A = 0; _arr_9260A <= 0; _arr_9260A = _arr_9260A + 1) begin : core_bus2_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_9260A_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_9260A_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [178:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [130:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache.sv:56:5
											wire [0:0] per_bank_flush_begin;
											// Trace: src/VX_cache.sv:57:5
											wire [0:0] flush_uuid;
											// Trace: src/VX_cache.sv:58:5
											wire [0:0] per_bank_flush_end;
											// Trace: src/VX_cache.sv:59:5
											wire [0:0] per_bank_core_req_fire;
											// Trace: src/VX_cache.sv:60:5
											// expanded module instance: flush_unit
											localparam _bbase_1DACF_core_bus_in_if = 0;
											localparam _bbase_1DACF_core_bus_out_if = 0;
											localparam _param_1DACF_NUM_REQS = NUM_REQS;
											localparam _param_1DACF_NUM_BANKS = NUM_BANKS;
											localparam _param_1DACF_UUID_WIDTH = UUID_WIDTH;
											localparam _param_1DACF_TAG_WIDTH = TAG_WIDTH;
											localparam _param_1DACF_BANK_SEL_LATENCY = 0;
											if (1) begin : flush_unit
												// Trace: src/VX_cache_flush.sv:2:15
												localparam NUM_REQS = _param_1DACF_NUM_REQS;
												// Trace: src/VX_cache_flush.sv:3:15
												localparam NUM_BANKS = _param_1DACF_NUM_BANKS;
												// Trace: src/VX_cache_flush.sv:4:15
												localparam UUID_WIDTH = _param_1DACF_UUID_WIDTH;
												// Trace: src/VX_cache_flush.sv:5:15
												localparam TAG_WIDTH = _param_1DACF_TAG_WIDTH;
												// Trace: src/VX_cache_flush.sv:6:15
												localparam BANK_SEL_LATENCY = _param_1DACF_BANK_SEL_LATENCY;
												// Trace: src/VX_cache_flush.sv:8:5
												wire clk;
												// Trace: src/VX_cache_flush.sv:9:5
												wire reset;
												// Trace: src/VX_cache_flush.sv:10:5
												localparam _mbase_core_bus_in_if = 0;
												// Trace: src/VX_cache_flush.sv:11:5
												localparam _mbase_core_bus_out_if = 0;
												// Trace: src/VX_cache_flush.sv:12:5
												wire [0:0] bank_req_fire;
												// Trace: src/VX_cache_flush.sv:13:5
												wire [0:0] flush_begin;
												// Trace: src/VX_cache_flush.sv:14:5
												wire [0:0] flush_uuid;
												// Trace: src/VX_cache_flush.sv:15:5
												wire [0:0] flush_end;
												// Trace: src/VX_cache_flush.sv:17:5
												localparam STATE_IDLE = 0;
												// Trace: src/VX_cache_flush.sv:18:5
												localparam STATE_WAIT1 = 1;
												// Trace: src/VX_cache_flush.sv:19:5
												localparam STATE_FLUSH = 2;
												// Trace: src/VX_cache_flush.sv:20:5
												localparam STATE_WAIT2 = 3;
												// Trace: src/VX_cache_flush.sv:21:5
												localparam STATE_DONE = 4;
												// Trace: src/VX_cache_flush.sv:22:5
												reg [2:0] state;
												reg [2:0] state_n;
												// Trace: src/VX_cache_flush.sv:23:5
												wire no_inflight_reqs;
												// Trace: src/VX_cache_flush.sv:24:5
												if (1) begin : g_no_bank_sel_latency
													// Trace: src/VX_cache_flush.sv:63:9
													assign no_inflight_reqs = 0;
												end
												// Trace: src/VX_cache_flush.sv:65:5
												reg [0:0] flush_done;
												reg [0:0] flush_done_n;
												// Trace: src/VX_cache_flush.sv:66:5
												wire [0:0] flush_req_mask;
												// Trace: src/VX_cache_flush.sv:67:5
												genvar _gv_i_116;
												for (_gv_i_116 = 0; _gv_i_116 < NUM_REQS; _gv_i_116 = _gv_i_116 + 1) begin : g_flush_req_mask
													localparam i = _gv_i_116;
													// Trace: src/VX_cache_flush.sv:68:9
													assign flush_req_mask[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data[3];
												end
												// Trace: src/VX_cache_flush.sv:70:5
												wire flush_req_enable = |flush_req_mask;
												// Trace: src/VX_cache_flush.sv:71:5
												reg [0:0] lock_released;
												reg [0:0] lock_released_n;
												// Trace: src/VX_cache_flush.sv:72:5
												reg [0:0] flush_uuid_r;
												reg [0:0] flush_uuid_n;
												// Trace: src/VX_cache_flush.sv:73:5
												genvar _gv_i_117;
												for (_gv_i_117 = 0; _gv_i_117 < NUM_REQS; _gv_i_117 = _gv_i_117 + 1) begin : g_core_bus_out_req
													localparam i = _gv_i_117;
													// Trace: src/VX_cache_flush.sv:74:9
													wire input_enable = ~flush_req_enable || lock_released[i];
													// Trace: src/VX_cache_flush.sv:75:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_valid && input_enable;
													// Trace: src/VX_cache_flush.sv:76:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data;
													// Trace: src/VX_cache_flush.sv:77:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_ready && input_enable;
												end
												// Trace: src/VX_cache_flush.sv:79:5
												genvar _gv_i_118;
												for (_gv_i_118 = 0; _gv_i_118 < NUM_REQS; _gv_i_118 = _gv_i_118 + 1) begin : g_core_bus_in_rsp
													localparam i = _gv_i_118;
													// Trace: src/VX_cache_flush.sv:80:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_valid;
													// Trace: src/VX_cache_flush.sv:81:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_data;
													// Trace: src/VX_cache_flush.sv:82:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_ready;
												end
												// Trace: src/VX_cache_flush.sv:84:5
												reg [0:0] core_bus_out_uuid;
												// Trace: src/VX_cache_flush.sv:85:5
												wire [0:0] core_bus_out_ready;
												// Trace: src/VX_cache_flush.sv:86:5
												genvar _gv_i_119;
												for (_gv_i_119 = 0; _gv_i_119 < NUM_REQS; _gv_i_119 = _gv_i_119 + 1) begin : g_core_bus_out_uuid
													localparam i = _gv_i_119;
													if (1) begin : g_uuid
														// Trace: src/VX_cache_flush.sv:88:13
														wire [1:1] sv2v_tmp_284C0;
														assign sv2v_tmp_284C0 = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data[2-:1];
														always @(*) core_bus_out_uuid[i+:1] = sv2v_tmp_284C0;
													end
												end
												// Trace: src/VX_cache_flush.sv:93:5
												genvar _gv_i_120;
												for (_gv_i_120 = 0; _gv_i_120 < NUM_REQS; _gv_i_120 = _gv_i_120 + 1) begin : g_core_bus_out_ready
													localparam i = _gv_i_120;
													// Trace: src/VX_cache_flush.sv:94:9
													assign core_bus_out_ready[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_ready;
												end
												// Trace: src/VX_cache_flush.sv:96:5
												always @(*) begin
													// Trace: src/VX_cache_flush.sv:97:9
													state_n = state;
													// Trace: src/VX_cache_flush.sv:98:9
													flush_done_n = flush_done;
													// Trace: src/VX_cache_flush.sv:99:9
													lock_released_n = lock_released;
													// Trace: src/VX_cache_flush.sv:100:9
													flush_uuid_n = flush_uuid_r;
													// Trace: src/VX_cache_flush.sv:101:9
													case (state)
														default:
															// Trace: src/VX_cache_flush.sv:103:17
															if (flush_req_enable) begin
																// Trace: src/VX_cache_flush.sv:104:21
																state_n = STATE_FLUSH;
																// Trace: src/VX_cache_flush.sv:105:21
																begin : sv2v_autoblock_2
																	// Trace: src/VX_cache_flush.sv:105:26
																	integer i;
																	// Trace: src/VX_cache_flush.sv:105:26
																	for (i = 0; i >= 0; i = i - 1)
																		begin
																			// Trace: src/VX_cache_flush.sv:106:25
																			if (flush_req_mask[i])
																				// Trace: src/VX_cache_flush.sv:107:29
																				flush_uuid_n = core_bus_out_uuid[i+:1];
																		end
																end
															end
														STATE_WAIT1:
															// Trace: src/VX_cache_flush.sv:113:17
															if (no_inflight_reqs)
																// Trace: src/VX_cache_flush.sv:114:21
																state_n = STATE_FLUSH;
														STATE_FLUSH:
															// Trace: src/VX_cache_flush.sv:118:17
															state_n = STATE_WAIT2;
														STATE_WAIT2: begin
															// Trace: src/VX_cache_flush.sv:121:17
															flush_done_n = flush_done | flush_end;
															// Trace: src/VX_cache_flush.sv:122:17
															if (flush_done_n == {NUM_BANKS {1'b1}}) begin
																// Trace: src/VX_cache_flush.sv:123:21
																state_n = STATE_DONE;
																// Trace: src/VX_cache_flush.sv:124:21
																flush_done_n = 1'sb0;
																// Trace: src/VX_cache_flush.sv:125:21
																lock_released_n = flush_req_mask;
															end
														end
														STATE_DONE: begin
															// Trace: src/VX_cache_flush.sv:129:17
															lock_released_n = lock_released & ~core_bus_out_ready;
															// Trace: src/VX_cache_flush.sv:130:17
															if (lock_released_n == 0)
																// Trace: src/VX_cache_flush.sv:131:21
																state_n = STATE_IDLE;
														end
													endcase
												end
												// Trace: src/VX_cache_flush.sv:136:5
												always @(posedge clk) begin
													// Trace: src/VX_cache_flush.sv:137:9
													if (reset) begin
														// Trace: src/VX_cache_flush.sv:138:13
														state <= STATE_IDLE;
														// Trace: src/VX_cache_flush.sv:139:13
														flush_done <= 1'sb0;
														// Trace: src/VX_cache_flush.sv:140:13
														lock_released <= 1'sb0;
													end
													else begin
														// Trace: src/VX_cache_flush.sv:142:13
														state <= state_n;
														// Trace: src/VX_cache_flush.sv:143:13
														flush_done <= flush_done_n;
														// Trace: src/VX_cache_flush.sv:144:13
														lock_released <= lock_released_n;
													end
													// Trace: src/VX_cache_flush.sv:146:9
													flush_uuid_r <= flush_uuid_n;
												end
												// Trace: src/VX_cache_flush.sv:148:5
												assign flush_begin = {NUM_BANKS {state == STATE_FLUSH}};
												// Trace: src/VX_cache_flush.sv:149:5
												assign flush_uuid = flush_uuid_r;
											end
											assign flush_unit.clk = clk;
											assign flush_unit.reset = reset;
											assign flush_unit.bank_req_fire = per_bank_core_req_fire;
											assign per_bank_flush_begin = flush_unit.flush_begin;
											assign flush_uuid = flush_unit.flush_uuid;
											assign flush_unit.flush_end = per_bank_flush_end;
											// Trace: src/VX_cache.sv:76:5
											// expanded interface instance: mem_bus_tmp_if
											localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
											localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
											genvar _arr_4FE36;
											for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam FLAGS_WIDTH = 3;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:7:15
												localparam UUID_WIDTH = 1;
												// Trace: src/VX_mem_bus_if.sv:9:5
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:13:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:21:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire [610:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire [516:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:30:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:31:5
												// Trace: src/VX_mem_bus_if.sv:39:5
											end
											// Trace: src/VX_cache.sv:80:5
											wire [0:0] mem_rsp_queue_valid;
											// Trace: src/VX_cache.sv:81:5
											wire [516:0] mem_rsp_queue_data;
											// Trace: src/VX_cache.sv:82:5
											wire [0:0] mem_rsp_queue_ready;
											// Trace: src/VX_cache.sv:83:5
											genvar _gv_i_29;
											for (_gv_i_29 = 0; _gv_i_29 < MEM_PORTS; _gv_i_29 = _gv_i_29 + 1) begin : g_mem_rsp_queue
												localparam i = _gv_i_29;
												// Trace: src/VX_cache.sv:84:9
												VX_elastic_buffer #(
													.DATAW(MEM_RSP_DATAW),
													.SIZE(MRSQ_SIZE),
													.OUT_REG(1'd1)
												) mem_rsp_queue(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_bus_tmp_if[i].rsp_valid),
													.data_in(mem_bus_tmp_if[i].rsp_data),
													.ready_in(mem_bus_tmp_if[i].rsp_ready),
													.valid_out(mem_rsp_queue_valid[i]),
													.data_out(mem_rsp_queue_data[i * 517+:517]),
													.ready_out(mem_rsp_queue_ready[i])
												);
											end
											// Trace: src/VX_cache.sv:99:5
											wire [516:0] mem_rsp_queue_data_s;
											// Trace: src/VX_cache.sv:100:5
											wire [0:0] mem_rsp_queue_sel;
											// Trace: src/VX_cache.sv:101:5
											genvar _gv_i_30;
											for (_gv_i_30 = 0; _gv_i_30 < MEM_PORTS; _gv_i_30 = _gv_i_30 + 1) begin : g_mem_rsp_queue_data_s
												localparam i = _gv_i_30;
												// Trace: src/VX_cache.sv:102:9
												wire [4:0] mem_rsp_tag_s = mem_rsp_queue_data[(i * 517) + 4-:5];
												// Trace: src/VX_cache.sv:103:9
												wire [511:0] mem_rsp_data_s = mem_rsp_queue_data[(i * 517) + 516-:512];
												// Trace: src/VX_cache.sv:104:9
												assign mem_rsp_queue_data_s[i * 517+:517] = {mem_rsp_data_s, mem_rsp_tag_s};
											end
											// Trace: src/VX_cache.sv:106:5
											genvar _gv_i_31;
											for (_gv_i_31 = 0; _gv_i_31 < MEM_PORTS; _gv_i_31 = _gv_i_31 + 1) begin : g_mem_rsp_queue_sel
												localparam i = _gv_i_31;
												if (1) begin : g_singlebank
													// Trace: src/VX_cache.sv:121:13
													assign mem_rsp_queue_sel[i+:1] = 0;
												end
											end
											// Trace: src/VX_cache.sv:124:5
											wire [0:0] per_bank_mem_rsp_valid;
											// Trace: src/VX_cache.sv:125:5
											wire [516:0] per_bank_mem_rsp_pdata;
											// Trace: src/VX_cache.sv:126:5
											wire [0:0] per_bank_mem_rsp_ready;
											// Trace: src/VX_cache.sv:127:5
											VX_stream_omega #(
												.NUM_INPUTS(MEM_PORTS),
												.NUM_OUTPUTS(NUM_BANKS),
												.DATAW(517),
												.ARBITER("R"),
												.OUT_BUF(3)
											) mem_rsp_xbar(
												.clk(clk),
												.reset(reset),
												.valid_in(mem_rsp_queue_valid),
												.data_in(mem_rsp_queue_data_s),
												.sel_in(mem_rsp_queue_sel),
												.ready_in(mem_rsp_queue_ready),
												.valid_out(per_bank_mem_rsp_valid),
												.data_out(per_bank_mem_rsp_pdata),
												.sel_out(),
												.ready_out(per_bank_mem_rsp_ready),
												.collisions()
											);
											// Trace: src/VX_cache.sv:146:5
											wire [511:0] per_bank_mem_rsp_data;
											// Trace: src/VX_cache.sv:147:5
											wire [4:0] per_bank_mem_rsp_tag;
											// Trace: src/VX_cache.sv:148:5
											genvar _gv_i_32;
											for (_gv_i_32 = 0; _gv_i_32 < NUM_BANKS; _gv_i_32 = _gv_i_32 + 1) begin : g_per_bank_mem_rsp_data
												localparam i = _gv_i_32;
												// Trace: src/VX_cache.sv:149:9
												assign {per_bank_mem_rsp_data[i * 512+:512], per_bank_mem_rsp_tag[i * 5+:5]} = per_bank_mem_rsp_pdata[i * 517+:517];
											end
											// Trace: src/VX_cache.sv:154:5
											wire [0:0] per_bank_core_req_valid;
											// Trace: src/VX_cache.sv:155:5
											wire [25:0] per_bank_core_req_addr;
											// Trace: src/VX_cache.sv:156:5
											wire [0:0] per_bank_core_req_rw;
											// Trace: src/VX_cache.sv:157:5
											wire [1:0] per_bank_core_req_wsel;
											// Trace: src/VX_cache.sv:158:5
											wire [15:0] per_bank_core_req_byteen;
											// Trace: src/VX_cache.sv:159:5
											wire [127:0] per_bank_core_req_data;
											// Trace: src/VX_cache.sv:160:5
											wire [2:0] per_bank_core_req_tag;
											// Trace: src/VX_cache.sv:161:5
											wire [0:0] per_bank_core_req_idx;
											// Trace: src/VX_cache.sv:162:5
											wire [2:0] per_bank_core_req_flags;
											// Trace: src/VX_cache.sv:163:5
											wire [0:0] per_bank_core_req_ready;
											// Trace: src/VX_cache.sv:164:5
											wire [0:0] per_bank_core_rsp_valid;
											// Trace: src/VX_cache.sv:165:5
											wire [127:0] per_bank_core_rsp_data;
											// Trace: src/VX_cache.sv:166:5
											wire [2:0] per_bank_core_rsp_tag;
											// Trace: src/VX_cache.sv:167:5
											wire [0:0] per_bank_core_rsp_idx;
											// Trace: src/VX_cache.sv:168:5
											wire [0:0] per_bank_core_rsp_ready;
											// Trace: src/VX_cache.sv:169:5
											wire [0:0] per_bank_mem_req_valid;
											// Trace: src/VX_cache.sv:170:5
											wire [25:0] per_bank_mem_req_addr;
											// Trace: src/VX_cache.sv:171:5
											wire [0:0] per_bank_mem_req_rw;
											// Trace: src/VX_cache.sv:172:5
											wire [63:0] per_bank_mem_req_byteen;
											// Trace: src/VX_cache.sv:173:5
											wire [511:0] per_bank_mem_req_data;
											// Trace: src/VX_cache.sv:174:5
											wire [4:0] per_bank_mem_req_tag;
											// Trace: src/VX_cache.sv:175:5
											wire [2:0] per_bank_mem_req_flags;
											// Trace: src/VX_cache.sv:176:5
											wire [0:0] per_bank_mem_req_ready;
											// Trace: src/VX_cache.sv:177:5
											wire [0:0] core_req_valid;
											// Trace: src/VX_cache.sv:178:5
											wire [27:0] core_req_addr;
											// Trace: src/VX_cache.sv:179:5
											wire [0:0] core_req_rw;
											// Trace: src/VX_cache.sv:180:5
											wire [15:0] core_req_byteen;
											// Trace: src/VX_cache.sv:181:5
											wire [127:0] core_req_data;
											// Trace: src/VX_cache.sv:182:5
											wire [2:0] core_req_tag;
											// Trace: src/VX_cache.sv:183:5
											wire [2:0] core_req_flags;
											// Trace: src/VX_cache.sv:184:5
											wire [0:0] core_req_ready;
											// Trace: src/VX_cache.sv:185:5
											wire [25:0] core_req_line_addr;
											// Trace: src/VX_cache.sv:186:5
											wire [0:0] core_req_bid;
											// Trace: src/VX_cache.sv:187:5
											wire [1:0] core_req_wsel;
											// Trace: src/VX_cache.sv:188:5
											wire [178:0] core_req_data_in;
											// Trace: src/VX_cache.sv:189:5
											wire [178:0] core_req_data_out;
											// Trace: src/VX_cache.sv:190:5
											genvar _gv_i_33;
											for (_gv_i_33 = 0; _gv_i_33 < NUM_REQS; _gv_i_33 = _gv_i_33 + 1) begin : g_core_req
												localparam i = _gv_i_33;
												// Trace: src/VX_cache.sv:191:9
												assign core_req_valid[i] = core_bus2_if[i].req_valid;
												// Trace: src/VX_cache.sv:192:9
												assign core_req_rw[i] = core_bus2_if[i].req_data[178];
												// Trace: src/VX_cache.sv:193:9
												assign core_req_byteen[i * 16+:16] = core_bus2_if[i].req_data[21-:16];
												// Trace: src/VX_cache.sv:194:9
												assign core_req_addr[i * 28+:28] = core_bus2_if[i].req_data[177-:28];
												// Trace: src/VX_cache.sv:195:9
												assign core_req_data[i * 128+:128] = core_bus2_if[i].req_data[149-:128];
												// Trace: src/VX_cache.sv:196:9
												assign core_req_tag[i * 3+:3] = core_bus2_if[i].req_data[2-:3];
												// Trace: src/VX_cache.sv:197:9
												assign core_req_flags[i * 3+:3] = sv2v_cast_3(core_bus2_if[i].req_data[5-:3]);
												// Trace: src/VX_cache.sv:198:9
												assign core_bus2_if[i].req_ready = core_req_ready[i];
											end
											// Trace: src/VX_cache.sv:200:5
											genvar _gv_i_34;
											for (_gv_i_34 = 0; _gv_i_34 < NUM_REQS; _gv_i_34 = _gv_i_34 + 1) begin : g_core_req_wsel
												localparam i = _gv_i_34;
												if (1) begin : g_wsel
													// Trace: src/VX_cache.sv:202:13
													assign core_req_wsel[i * 2+:2] = core_req_addr[i * 28+:WORD_SEL_BITS];
												end
											end
											// Trace: src/VX_cache.sv:207:5
											genvar _gv_i_35;
											for (_gv_i_35 = 0; _gv_i_35 < NUM_REQS; _gv_i_35 = _gv_i_35 + 1) begin : g_core_req_line_addr
												localparam i = _gv_i_35;
												// Trace: src/VX_cache.sv:208:9
												assign core_req_line_addr[i * 26+:26] = core_req_addr[(i * 28) + 2+:LINE_ADDR_WIDTH];
											end
											// Trace: src/VX_cache.sv:210:5
											genvar _gv_i_36;
											for (_gv_i_36 = 0; _gv_i_36 < NUM_REQS; _gv_i_36 = _gv_i_36 + 1) begin : g_core_req_bid
												localparam i = _gv_i_36;
												if (1) begin : g_singlebank
													// Trace: src/VX_cache.sv:214:13
													assign core_req_bid[i+:1] = 1'sb0;
												end
											end
											// Trace: src/VX_cache.sv:217:5
											genvar _gv_i_37;
											for (_gv_i_37 = 0; _gv_i_37 < NUM_REQS; _gv_i_37 = _gv_i_37 + 1) begin : g_core_req_data_in
												localparam i = _gv_i_37;
												// Trace: src/VX_cache.sv:218:9
												assign core_req_data_in[i * 179+:179] = {core_req_line_addr[i * 26+:26], core_req_rw[i], core_req_wsel[i * 2+:2], core_req_byteen[i * 16+:16], core_req_data[i * 128+:128], core_req_tag[i * 3+:3], core_req_flags[i * 3+:3]};
											end
											// Trace: src/VX_cache.sv:228:5
											assign per_bank_core_req_fire = per_bank_core_req_valid & per_bank_mem_req_ready;
											// Trace: src/VX_cache.sv:229:5
											VX_stream_xbar #(
												.NUM_INPUTS(NUM_REQS),
												.NUM_OUTPUTS(NUM_BANKS),
												.DATAW(CORE_REQ_DATAW),
												.PERF_CTR_BITS(44),
												.ARBITER("R"),
												.OUT_BUF(REQ_XBAR_BUF)
											) req_xbar(
												.clk(clk),
												.reset(reset),
												.collisions(),
												.valid_in(core_req_valid),
												.data_in(core_req_data_in),
												.sel_in(core_req_bid),
												.ready_in(core_req_ready),
												.valid_out(per_bank_core_req_valid),
												.data_out(core_req_data_out),
												.sel_out(per_bank_core_req_idx),
												.ready_out(per_bank_core_req_ready)
											);
											// Trace: src/VX_cache.sv:249:5
											genvar _gv_i_38;
											for (_gv_i_38 = 0; _gv_i_38 < NUM_BANKS; _gv_i_38 = _gv_i_38 + 1) begin : g_core_req_data_out
												localparam i = _gv_i_38;
												// Trace: src/VX_cache.sv:250:9
												assign {per_bank_core_req_addr[i * 26+:26], per_bank_core_req_rw[i], per_bank_core_req_wsel[i * 2+:2], per_bank_core_req_byteen[i * 16+:16], per_bank_core_req_data[i * 128+:128], per_bank_core_req_tag[i * 3+:3], per_bank_core_req_flags[i * 3+:3]} = core_req_data_out[i * 179+:179];
											end
											// Trace: src/VX_cache.sv:260:5
											genvar _gv_bank_id_1;
											for (_gv_bank_id_1 = 0; _gv_bank_id_1 < NUM_BANKS; _gv_bank_id_1 = _gv_bank_id_1 + 1) begin : g_banks
												localparam bank_id = _gv_bank_id_1;
												// Trace: src/VX_cache.sv:261:9
												VX_cache_bank #(
													.BANK_ID(bank_id),
													.INSTANCE_ID(""),
													.CACHE_SIZE(CACHE_SIZE),
													.LINE_SIZE(LINE_SIZE),
													.NUM_BANKS(NUM_BANKS),
													.NUM_WAYS(NUM_WAYS),
													.WORD_SIZE(WORD_SIZE),
													.NUM_REQS(NUM_REQS),
													.WRITE_ENABLE(WRITE_ENABLE),
													.WRITEBACK(WRITEBACK),
													.DIRTY_BYTES(DIRTY_BYTES),
													.REPL_POLICY(REPL_POLICY),
													.CRSQ_SIZE(CRSQ_SIZE),
													.MSHR_SIZE(MSHR_SIZE),
													.MREQ_SIZE(MREQ_SIZE),
													.UUID_WIDTH(UUID_WIDTH),
													.TAG_WIDTH(TAG_WIDTH),
													.FLAGS_WIDTH(FLAGS_WIDTH),
													.CORE_OUT_REG((CORE_RSP_REG_DISABLE ? 0 : 1)),
													.MEM_OUT_REG((MEM_REQ_REG_DISABLE ? 0 : 1))
												) bank(
													.clk(clk),
													.reset(reset),
													.core_req_valid(per_bank_core_req_valid[bank_id]),
													.core_req_addr(per_bank_core_req_addr[bank_id * 26+:26]),
													.core_req_rw(per_bank_core_req_rw[bank_id]),
													.core_req_wsel(per_bank_core_req_wsel[bank_id * 2+:2]),
													.core_req_byteen(per_bank_core_req_byteen[bank_id * 16+:16]),
													.core_req_data(per_bank_core_req_data[bank_id * 128+:128]),
													.core_req_tag(per_bank_core_req_tag[bank_id * 3+:3]),
													.core_req_idx(per_bank_core_req_idx[bank_id+:1]),
													.core_req_flags(per_bank_core_req_flags[bank_id * 3+:3]),
													.core_req_ready(per_bank_core_req_ready[bank_id]),
													.core_rsp_valid(per_bank_core_rsp_valid[bank_id]),
													.core_rsp_data(per_bank_core_rsp_data[bank_id * 128+:128]),
													.core_rsp_tag(per_bank_core_rsp_tag[bank_id * 3+:3]),
													.core_rsp_idx(per_bank_core_rsp_idx[bank_id+:1]),
													.core_rsp_ready(per_bank_core_rsp_ready[bank_id]),
													.mem_req_valid(per_bank_mem_req_valid[bank_id]),
													.mem_req_addr(per_bank_mem_req_addr[bank_id * 26+:26]),
													.mem_req_rw(per_bank_mem_req_rw[bank_id]),
													.mem_req_byteen(per_bank_mem_req_byteen[bank_id * 64+:64]),
													.mem_req_data(per_bank_mem_req_data[bank_id * 512+:512]),
													.mem_req_tag(per_bank_mem_req_tag[bank_id * 5+:5]),
													.mem_req_flags(per_bank_mem_req_flags[bank_id * 3+:3]),
													.mem_req_ready(per_bank_mem_req_ready[bank_id]),
													.mem_rsp_valid(per_bank_mem_rsp_valid[bank_id]),
													.mem_rsp_data(per_bank_mem_rsp_data[bank_id * 512+:512]),
													.mem_rsp_tag(per_bank_mem_rsp_tag[bank_id * 5+:5]),
													.mem_rsp_ready(per_bank_mem_rsp_ready[bank_id]),
													.flush_begin(per_bank_flush_begin[bank_id]),
													.flush_uuid(flush_uuid),
													.flush_end(per_bank_flush_end[bank_id])
												);
											end
											// Trace: src/VX_cache.sv:317:5
											wire [130:0] core_rsp_data_in;
											// Trace: src/VX_cache.sv:318:5
											wire [130:0] core_rsp_data_out;
											// Trace: src/VX_cache.sv:319:5
											wire [0:0] core_rsp_valid_s;
											// Trace: src/VX_cache.sv:320:5
											wire [127:0] core_rsp_data_s;
											// Trace: src/VX_cache.sv:321:5
											wire [2:0] core_rsp_tag_s;
											// Trace: src/VX_cache.sv:322:5
											wire [0:0] core_rsp_ready_s;
											// Trace: src/VX_cache.sv:323:5
											genvar _gv_i_39;
											for (_gv_i_39 = 0; _gv_i_39 < NUM_BANKS; _gv_i_39 = _gv_i_39 + 1) begin : g_core_rsp_data_in
												localparam i = _gv_i_39;
												// Trace: src/VX_cache.sv:324:9
												assign core_rsp_data_in[i * 131+:131] = {per_bank_core_rsp_data[i * 128+:128], per_bank_core_rsp_tag[i * 3+:3]};
											end
											// Trace: src/VX_cache.sv:326:5
											VX_stream_xbar #(
												.NUM_INPUTS(NUM_BANKS),
												.NUM_OUTPUTS(NUM_REQS),
												.DATAW(CORE_RSP_DATAW),
												.ARBITER("R")
											) rsp_xbar(
												.clk(clk),
												.reset(reset),
												.collisions(),
												.valid_in(per_bank_core_rsp_valid),
												.data_in(core_rsp_data_in),
												.sel_in(per_bank_core_rsp_idx),
												.ready_in(per_bank_core_rsp_ready),
												.valid_out(core_rsp_valid_s),
												.data_out(core_rsp_data_out),
												.ready_out(core_rsp_ready_s),
												.sel_out()
											);
											// Trace: src/VX_cache.sv:344:5
											genvar _gv_i_40;
											for (_gv_i_40 = 0; _gv_i_40 < NUM_REQS; _gv_i_40 = _gv_i_40 + 1) begin : g_core_rsp_data_s
												localparam i = _gv_i_40;
												// Trace: src/VX_cache.sv:345:9
												assign {core_rsp_data_s[i * 128+:128], core_rsp_tag_s[i * 3+:3]} = core_rsp_data_out[i * 131+:131];
											end
											// Trace: src/VX_cache.sv:347:5
											genvar _gv_i_41;
											for (_gv_i_41 = 0; _gv_i_41 < NUM_REQS; _gv_i_41 = _gv_i_41 + 1) begin : g_core_rsp_buf
												localparam i = _gv_i_41;
												// Trace: src/VX_cache.sv:348:9
												VX_elastic_buffer #(
													.DATAW(131),
													.SIZE((CORE_RSP_REG_DISABLE ? ((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : 2) : 0)),
													.OUT_REG(((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : (CORE_OUT_BUF & 7) - 2))
												) core_rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(core_rsp_valid_s[i]),
													.ready_in(core_rsp_ready_s[i]),
													.data_in({core_rsp_data_s[i * 128+:128], core_rsp_tag_s[i * 3+:3]}),
													.data_out({core_bus2_if[i].rsp_data[130-:128], core_bus2_if[i].rsp_data[2-:3]}),
													.valid_out(core_bus2_if[i].rsp_valid),
													.ready_out(core_bus2_if[i].rsp_ready)
												);
											end
											// Trace: src/VX_cache.sv:363:5
											wire [610:0] per_bank_mem_req_pdata;
											// Trace: src/VX_cache.sv:364:5
											genvar _gv_i_42;
											for (_gv_i_42 = 0; _gv_i_42 < NUM_BANKS; _gv_i_42 = _gv_i_42 + 1) begin : g_per_bank_mem_req_pdata
												localparam i = _gv_i_42;
												// Trace: src/VX_cache.sv:365:9
												assign per_bank_mem_req_pdata[i * 611+:611] = {per_bank_mem_req_rw[i], per_bank_mem_req_addr[i * 26+:26], per_bank_mem_req_data[i * 512+:512], per_bank_mem_req_byteen[i * 64+:64], per_bank_mem_req_flags[i * 3+:3], per_bank_mem_req_tag[i * 5+:5]};
											end
											// Trace: src/VX_cache.sv:374:5
											wire [0:0] mem_req_valid;
											// Trace: src/VX_cache.sv:375:5
											wire [610:0] mem_req_pdata;
											// Trace: src/VX_cache.sv:376:5
											wire [0:0] mem_req_ready;
											// Trace: src/VX_cache.sv:377:5
											wire [0:0] mem_req_sel_out;
											// Trace: src/VX_cache.sv:378:5
											VX_stream_arb #(
												.NUM_INPUTS(NUM_BANKS),
												.NUM_OUTPUTS(MEM_PORTS),
												.DATAW(MEM_REQ_DATAW),
												.ARBITER("R")
											) mem_req_arb(
												.clk(clk),
												.reset(reset),
												.valid_in(per_bank_mem_req_valid),
												.data_in(per_bank_mem_req_pdata),
												.ready_in(per_bank_mem_req_ready),
												.valid_out(mem_req_valid),
												.data_out(mem_req_pdata),
												.ready_out(mem_req_ready),
												.sel_out(mem_req_sel_out)
											);
											// Trace: src/VX_cache.sv:394:5
											genvar _gv_i_43;
											for (_gv_i_43 = 0; _gv_i_43 < MEM_PORTS; _gv_i_43 = _gv_i_43 + 1) begin : g_mem_req_buf
												localparam i = _gv_i_43;
												// Trace: src/VX_cache.sv:395:9
												wire mem_req_rw;
												// Trace: src/VX_cache.sv:396:9
												wire [25:0] mem_req_addr;
												// Trace: src/VX_cache.sv:397:9
												wire [511:0] mem_req_data;
												// Trace: src/VX_cache.sv:398:9
												wire [63:0] mem_req_byteen;
												// Trace: src/VX_cache.sv:399:9
												wire [2:0] mem_req_flags;
												// Trace: src/VX_cache.sv:400:9
												wire [4:0] mem_req_tag;
												// Trace: src/VX_cache.sv:401:9
												assign {mem_req_rw, mem_req_addr, mem_req_data, mem_req_byteen, mem_req_flags, mem_req_tag} = mem_req_pdata[i * 611+:611];
												// Trace: src/VX_cache.sv:409:9
												wire [25:0] mem_req_addr_w;
												// Trace: src/VX_cache.sv:410:9
												wire [4:0] mem_req_tag_w;
												// Trace: src/VX_cache.sv:411:9
												wire [2:0] mem_req_flags_w;
												if (1) begin : g_mem_req_tag
													// Trace: src/VX_cache.sv:430:13
													assign mem_req_addr_w = mem_req_addr;
													// Trace: src/VX_cache.sv:431:13
													assign mem_req_tag_w = mem_req_tag;
												end
												// Trace: src/VX_cache.sv:433:9
												VX_elastic_buffer #(
													.DATAW(611),
													.SIZE((MEM_REQ_REG_DISABLE ? ((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : 2) : 0)),
													.OUT_REG(((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : (MEM_OUT_BUF & 7) - 2))
												) mem_req_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_req_valid[i]),
													.ready_in(mem_req_ready[i]),
													.data_in({mem_req_rw, mem_req_byteen, mem_req_addr_w, mem_req_data, mem_req_tag_w, mem_req_flags}),
													.data_out({mem_bus_tmp_if[i].req_data[610], mem_bus_tmp_if[i].req_data[71-:64], mem_bus_tmp_if[i].req_data[609-:26], mem_bus_tmp_if[i].req_data[583-:512], mem_bus_tmp_if[i].req_data[4-:5], mem_req_flags_w}),
													.valid_out(mem_bus_tmp_if[i].req_valid),
													.ready_out(mem_bus_tmp_if[i].req_ready)
												);
												if (1) begin : g_mem_req_flags
													// Trace: src/VX_cache.sv:448:13
													assign mem_bus_tmp_if[i].req_data[7-:3] = mem_req_flags_w;
												end
												if (WRITE_ENABLE) begin : g_mem_bus_if
													// Trace: src/VX_cache.sv:453:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
													// Trace: src/VX_cache.sv:454:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
													// Trace: src/VX_cache.sv:455:5
													assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_ready;
													// Trace: src/VX_cache.sv:456:5
													assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_valid;
													// Trace: src/VX_cache.sv:457:5
													assign mem_bus_tmp_if[i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data;
													// Trace: src/VX_cache.sv:458:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
												end
												else begin : g_mem_bus_if_ro
													// Trace: src/VX_cache.sv:460:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
													// Trace: src/VX_cache.sv:461:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[610] = 0;
													// Trace: src/VX_cache.sv:462:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[609-:26] = mem_bus_tmp_if[i].req_data[609-:26];
													// Trace: src/VX_cache.sv:463:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[583-:512] = 1'sb0;
													// Trace: src/VX_cache.sv:464:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[71-:64] = 1'sb1;
													// Trace: src/VX_cache.sv:465:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[7-:3] = mem_bus_tmp_if[i].req_data[7-:3];
													// Trace: src/VX_cache.sv:466:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[4-:5] = mem_bus_tmp_if[i].req_data[4-:5];
													// Trace: src/VX_cache.sv:467:5
													assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_ready;
													// Trace: src/VX_cache.sv:468:5
													assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_valid;
													// Trace: src/VX_cache.sv:469:5
													assign mem_bus_tmp_if[i].rsp_data[516-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data[516-:512];
													// Trace: src/VX_cache.sv:470:5
													assign mem_bus_tmp_if[i].rsp_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data[4-:5];
													// Trace: src/VX_cache.sv:471:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_66].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
												end
											end
										end
										assign cache.clk = clk;
										assign cache.reset = reset;
									end
								end
								assign cache_wrap.clk = clk;
								assign cache_wrap.reset = reset;
							end
							// Trace: src/VX_cache_cluster.sv:124:5
							genvar _gv_i_67;
							for (_gv_i_67 = 0; _gv_i_67 < MEM_PORTS; _gv_i_67 = _gv_i_67 + 1) begin : g_mem_bus_if
								localparam i = _gv_i_67;
								// Trace: src/VX_cache_cluster.sv:125:9
								// expanded interface instance: arb_core_bus_tmp_if
								localparam _param_E788B_DATA_SIZE = LINE_SIZE;
								localparam _param_E788B_TAG_WIDTH = MEM_TAG_WIDTH;
								genvar _arr_E788B;
								for (_arr_E788B = 0; _arr_E788B <= 0; _arr_E788B = _arr_E788B + 1) begin : arb_core_bus_tmp_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_E788B_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_E788B_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [611:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [517:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								// Trace: src/VX_cache_cluster.sv:129:9
								// expanded interface instance: mem_bus_tmp_if
								localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
								localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH + 0;
								genvar _arr_4FE36;
								for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [611:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [517:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								genvar _gv_j_7;
								for (_gv_j_7 = 0; _gv_j_7 < NUM_CACHES; _gv_j_7 = _gv_j_7 + 1) begin : g_arb_core_bus_tmp_if
									localparam j = _gv_j_7;
									// Trace: src/VX_cache_cluster.sv:134:5
									assign arb_core_bus_tmp_if[j].req_valid = cache_mem_bus_if[(j * MEM_PORTS) + i].req_valid;
									// Trace: src/VX_cache_cluster.sv:135:5
									assign arb_core_bus_tmp_if[j].req_data = cache_mem_bus_if[(j * MEM_PORTS) + i].req_data;
									// Trace: src/VX_cache_cluster.sv:136:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].req_ready = arb_core_bus_tmp_if[j].req_ready;
									// Trace: src/VX_cache_cluster.sv:137:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_valid = arb_core_bus_tmp_if[j].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:138:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_data = arb_core_bus_tmp_if[j].rsp_data;
									// Trace: src/VX_cache_cluster.sv:139:5
									assign arb_core_bus_tmp_if[j].rsp_ready = cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_ready;
								end
								// Trace: src/VX_cache_cluster.sv:141:9
								// expanded module instance: mem_arb
								localparam _bbase_7277A_bus_in_if = 0;
								localparam _bbase_7277A_bus_out_if = 0;
								localparam _param_7277A_NUM_INPUTS = NUM_CACHES;
								localparam _param_7277A_NUM_OUTPUTS = 1;
								localparam _param_7277A_DATA_SIZE = LINE_SIZE;
								localparam _param_7277A_TAG_WIDTH = MEM_TAG_WIDTH;
								localparam _param_7277A_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_7277A_ARBITER = "R";
								localparam _param_7277A_REQ_OUT_BUF = 0;
								localparam _param_7277A_RSP_OUT_BUF = 0;
								if (1) begin : mem_arb
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_7277A_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = _param_7277A_NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_7277A_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_7277A_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_7277A_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_7277A_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_7277A_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:16
									localparam ARBITER = _param_7277A_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 512;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 0;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 606 + TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [0:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [REQ_DATAW - 1:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [0:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [REQ_DATAW - 1:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_80;
									for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
										localparam i = _gv_i_80;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 612+:612] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_81;
									for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
										localparam i = _gv_i_81;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [TAG_WIDTH - 1:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										VX_bits_insert #(
											.N(TAG_WIDTH),
											.S(LOG_NUM_REQS),
											.POS(TAG_SEL_IDX)
										) bits_insert(
											.data_in(req_tag_out),
											.ins_in(req_sel_out[i+:1]),
											.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[5-:6])
										);
										// Trace: src/VX_mem_arb.sv:64:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:65:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[611], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[610-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[584-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[72-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[8-:3], req_tag_out} = req_data_out[i * 612+:612];
										// Trace: src/VX_mem_arb.sv:73:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
									end
									// Trace: src/VX_mem_arb.sv:75:5
									wire [0:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:76:5
									wire [RSP_DATAW - 1:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:77:5
									wire [0:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:78:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:79:5
									wire [RSP_DATAW - 1:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:81:5
									if (1) begin : g_passthru
										genvar _gv_i_83;
										for (_gv_i_83 = 0; _gv_i_83 < NUM_OUTPUTS; _gv_i_83 = _gv_i_83 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_83;
											// Trace: src/VX_mem_arb.sv:116:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:117:13
											assign rsp_data_in[i * 518+:518] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
											// Trace: src/VX_mem_arb.sv:118:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:120:9
										VX_stream_arb #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.ARBITER(ARBITER),
											.OUT_BUF(RSP_OUT_BUF)
										) req_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
									end
									// Trace: src/VX_mem_arb.sv:138:5
									genvar _gv_i_84;
									for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
										localparam i = _gv_i_84;
										// Trace: src/VX_mem_arb.sv:139:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:140:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 518+:518];
										// Trace: src/VX_mem_arb.sv:141:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_67].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign mem_arb.clk = clk;
								assign mem_arb.reset = reset;
								if (WRITE_ENABLE) begin : g_we
									// Trace: src/VX_cache_cluster.sv:157:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[0].req_valid;
									// Trace: src/VX_cache_cluster.sv:158:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[0].req_data;
									// Trace: src/VX_cache_cluster.sv:159:5
									assign mem_bus_tmp_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
									// Trace: src/VX_cache_cluster.sv:160:5
									assign mem_bus_tmp_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:161:5
									assign mem_bus_tmp_if[0].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
									// Trace: src/VX_cache_cluster.sv:162:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[0].rsp_ready;
								end
								else begin : g_ro
									// Trace: src/VX_cache_cluster.sv:164:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[0].req_valid;
									// Trace: src/VX_cache_cluster.sv:165:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[611] = 0;
									// Trace: src/VX_cache_cluster.sv:166:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[610-:26] = mem_bus_tmp_if[0].req_data[610-:26];
									// Trace: src/VX_cache_cluster.sv:167:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[584-:512] = 1'sb0;
									// Trace: src/VX_cache_cluster.sv:168:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[72-:64] = 1'sb1;
									// Trace: src/VX_cache_cluster.sv:169:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[8-:3] = mem_bus_tmp_if[0].req_data[8-:3];
									// Trace: src/VX_cache_cluster.sv:170:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[5-:6] = mem_bus_tmp_if[0].req_data[5-:6];
									// Trace: src/VX_cache_cluster.sv:171:5
									assign mem_bus_tmp_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
									// Trace: src/VX_cache_cluster.sv:172:5
									assign mem_bus_tmp_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:173:5
									assign mem_bus_tmp_if[0].rsp_data[517-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[517-:512];
									// Trace: src/VX_cache_cluster.sv:174:5
									assign mem_bus_tmp_if[0].rsp_data[5-:6] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[5-:6];
									// Trace: src/VX_cache_cluster.sv:175:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[0].rsp_ready;
								end
							end
						end
						assign dcache.clk = clk;
						assign dcache.reset = dcache_reset;
						// Trace: src/VX_socket.sv:101:5
						genvar _gv_i_153;
						localparam VX_gpu_pkg_L1_MEM_TAG_WIDTH = VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH;
						localparam VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH = 7;
						for (_gv_i_153 = 0; _gv_i_153 < VX_gpu_pkg_DCACHE_NUM_REQS; _gv_i_153 = _gv_i_153 + 1) begin : g_mem_bus_if
							localparam i = _gv_i_153;
							if (i == 0) begin : g_i0
								// Trace: src/VX_socket.sv:103:13
								// expanded interface instance: l1_mem_bus_if
								localparam _param_70CB9_DATA_SIZE = 64;
								localparam _param_70CB9_TAG_WIDTH = VX_gpu_pkg_L1_MEM_TAG_WIDTH;
								genvar _arr_70CB9;
								for (_arr_70CB9 = 0; _arr_70CB9 <= 1; _arr_70CB9 = _arr_70CB9 + 1) begin : l1_mem_bus_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_70CB9_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_70CB9_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [611:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [517:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								// Trace: src/VX_socket.sv:107:13
								// expanded interface instance: l1_mem_arb_bus_if
								localparam _param_D5D25_DATA_SIZE = 64;
								localparam _param_D5D25_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
								genvar _arr_D5D25;
								for (_arr_D5D25 = 0; _arr_D5D25 <= 0; _arr_D5D25 = _arr_D5D25 + 1) begin : l1_mem_arb_bus_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_D5D25_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_D5D25_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [612:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [518:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								// Trace: src/VX_socket.sv:111:5
								assign l1_mem_bus_if[0].req_valid = icache_mem_bus_if[0].req_valid;
								// Trace: src/VX_socket.sv:112:5
								assign l1_mem_bus_if[0].req_data[611] = icache_mem_bus_if[0].req_data[610];
								// Trace: src/VX_socket.sv:113:5
								assign l1_mem_bus_if[0].req_data[610-:26] = icache_mem_bus_if[0].req_data[609-:26];
								// Trace: src/VX_socket.sv:114:5
								assign l1_mem_bus_if[0].req_data[584-:512] = icache_mem_bus_if[0].req_data[583-:512];
								// Trace: src/VX_socket.sv:115:5
								assign l1_mem_bus_if[0].req_data[72-:64] = icache_mem_bus_if[0].req_data[71-:64];
								// Trace: src/VX_socket.sv:116:5
								assign l1_mem_bus_if[0].req_data[8-:3] = icache_mem_bus_if[0].req_data[7-:3];
								if (1) begin : genblk1
									if (1) begin : genblk1
										if (1) begin : genblk1
											// Trace: src/VX_socket.sv:121:17
											assign l1_mem_bus_if[0].req_data[5-:6] = {icache_mem_bus_if[0].req_data[4-:1], 1'b0, icache_mem_bus_if[0].req_data[3-:4]};
										end
									end
								end
								// Trace: src/VX_socket.sv:136:5
								assign icache_mem_bus_if[0].req_ready = l1_mem_bus_if[0].req_ready;
								// Trace: src/VX_socket.sv:137:5
								assign icache_mem_bus_if[0].rsp_valid = l1_mem_bus_if[0].rsp_valid;
								// Trace: src/VX_socket.sv:138:5
								assign icache_mem_bus_if[0].rsp_data[516-:512] = l1_mem_bus_if[0].rsp_data[517-:512];
								if (1) begin : genblk2
									if (1) begin : genblk1
										if (1) begin : genblk1
											// Trace: src/VX_socket.sv:143:17
											assign icache_mem_bus_if[0].rsp_data[4-:5] = {l1_mem_bus_if[0].rsp_data[5-:1], l1_mem_bus_if[0].rsp_data[3:0]};
										end
									end
								end
								// Trace: src/VX_socket.sv:158:5
								assign l1_mem_bus_if[0].rsp_ready = icache_mem_bus_if[0].rsp_ready;
								// Trace: src/VX_socket.sv:159:5
								assign l1_mem_bus_if[1].req_valid = dcache_mem_bus_if[0].req_valid;
								// Trace: src/VX_socket.sv:160:5
								assign l1_mem_bus_if[1].req_data[611] = dcache_mem_bus_if[0].req_data[611];
								// Trace: src/VX_socket.sv:161:5
								assign l1_mem_bus_if[1].req_data[610-:26] = dcache_mem_bus_if[0].req_data[610-:26];
								// Trace: src/VX_socket.sv:162:5
								assign l1_mem_bus_if[1].req_data[584-:512] = dcache_mem_bus_if[0].req_data[584-:512];
								// Trace: src/VX_socket.sv:163:5
								assign l1_mem_bus_if[1].req_data[72-:64] = dcache_mem_bus_if[0].req_data[72-:64];
								// Trace: src/VX_socket.sv:164:5
								assign l1_mem_bus_if[1].req_data[8-:3] = dcache_mem_bus_if[0].req_data[8-:3];
								if (1) begin : genblk3
									// Trace: src/VX_socket.sv:181:9
									assign l1_mem_bus_if[1].req_data[5-:6] = dcache_mem_bus_if[0].req_data[5-:6];
								end
								// Trace: src/VX_socket.sv:184:5
								assign dcache_mem_bus_if[0].req_ready = l1_mem_bus_if[1].req_ready;
								// Trace: src/VX_socket.sv:185:5
								assign dcache_mem_bus_if[0].rsp_valid = l1_mem_bus_if[1].rsp_valid;
								// Trace: src/VX_socket.sv:186:5
								assign dcache_mem_bus_if[0].rsp_data[517-:512] = l1_mem_bus_if[1].rsp_data[517-:512];
								if (1) begin : genblk4
									// Trace: src/VX_socket.sv:203:9
									assign dcache_mem_bus_if[0].rsp_data[5-:6] = l1_mem_bus_if[1].rsp_data[5-:6];
								end
								// Trace: src/VX_socket.sv:206:5
								assign l1_mem_bus_if[1].rsp_ready = dcache_mem_bus_if[0].rsp_ready;
								// Trace: src/VX_socket.sv:207:13
								// expanded module instance: mem_arb
								localparam _bbase_7277A_bus_in_if = 0;
								localparam _bbase_7277A_bus_out_if = 0;
								localparam _param_7277A_NUM_INPUTS = 2;
								localparam _param_7277A_DATA_SIZE = 64;
								localparam _param_7277A_TAG_WIDTH = VX_gpu_pkg_L1_MEM_TAG_WIDTH;
								localparam _param_7277A_TAG_SEL_IDX = 0;
								localparam _param_7277A_ARBITER = "P";
								localparam _param_7277A_REQ_OUT_BUF = 3;
								localparam _param_7277A_RSP_OUT_BUF = 3;
								if (1) begin : mem_arb
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_7277A_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = 1;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_7277A_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_7277A_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_7277A_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_7277A_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_7277A_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:16
									localparam ARBITER = _param_7277A_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 512;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 1;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 612;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = 518;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [1:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [1223:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [1:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [611:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_80;
									for (_gv_i_80 = 0; _gv_i_80 < NUM_INPUTS; _gv_i_80 = _gv_i_80 + 1) begin : g_req_data_in
										localparam i = _gv_i_80;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 612+:612] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_81;
									for (_gv_i_81 = 0; _gv_i_81 < NUM_OUTPUTS; _gv_i_81 = _gv_i_81 + 1) begin : g_bus_out_if
										localparam i = _gv_i_81;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [5:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										VX_bits_insert #(
											.N(TAG_WIDTH),
											.S(LOG_NUM_REQS),
											.POS(TAG_SEL_IDX)
										) bits_insert(
											.data_in(req_tag_out),
											.ins_in(req_sel_out[i+:1]),
											.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[6-:7])
										);
										// Trace: src/VX_mem_arb.sv:64:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:65:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[612], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[611-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[585-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[73-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[9-:3], req_tag_out} = req_data_out[i * 612+:612];
										// Trace: src/VX_mem_arb.sv:73:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_ready;
									end
									// Trace: src/VX_mem_arb.sv:75:5
									wire [1:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:76:5
									wire [1035:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:77:5
									wire [1:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:78:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:79:5
									wire [517:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:81:5
									if (1) begin : g_rsp_enabled
										// Trace: src/VX_mem_arb.sv:82:9
										wire [0:0] rsp_sel_in;
										genvar _gv_i_82;
										for (_gv_i_82 = 0; _gv_i_82 < NUM_OUTPUTS; _gv_i_82 = _gv_i_82 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_82;
											// Trace: src/VX_mem_arb.sv:84:13
											wire [5:0] rsp_tag_out;
											// Trace: src/VX_mem_arb.sv:85:13
											VX_bits_remove #(
												.N(7),
												.S(LOG_NUM_REQS),
												.POS(TAG_SEL_IDX)
											) bits_remove(
												.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].rsp_data[6-:7]),
												.sel_out(rsp_sel_in[i+:1]),
												.data_out(rsp_tag_out)
											);
											// Trace: src/VX_mem_arb.sv:94:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:95:13
											assign rsp_data_in[i * 518+:518] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].rsp_data[518-:512], rsp_tag_out};
											// Trace: src/VX_mem_arb.sv:96:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:98:9
										VX_stream_switch #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.OUT_BUF(RSP_OUT_BUF)
										) rsp_switch(
											.clk(clk),
											.reset(reset),
											.sel_in(rsp_sel_in),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out)
										);
									end
									// Trace: src/VX_mem_arb.sv:138:5
									genvar _gv_i_84;
									for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_output
										localparam i = _gv_i_84;
										// Trace: src/VX_mem_arb.sv:139:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:140:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 518+:518];
										// Trace: src/VX_mem_arb.sv:141:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_153].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign mem_arb.clk = clk;
								assign mem_arb.reset = reset;
								// Trace: src/VX_socket.sv:221:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].req_valid = l1_mem_arb_bus_if[0].req_valid;
								// Trace: src/VX_socket.sv:222:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].req_data = l1_mem_arb_bus_if[0].req_data;
								// Trace: src/VX_socket.sv:223:5
								assign l1_mem_arb_bus_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].req_ready;
								// Trace: src/VX_socket.sv:224:5
								assign l1_mem_arb_bus_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].rsp_valid;
								// Trace: src/VX_socket.sv:225:5
								assign l1_mem_arb_bus_if[0].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].rsp_data;
								// Trace: src/VX_socket.sv:226:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].rsp_ready = l1_mem_arb_bus_if[0].rsp_ready;
							end
							else begin : g_i
								// Trace: src/VX_socket.sv:228:13
								// expanded interface instance: l1_mem_arb_bus_if
								localparam _param_D5D25_DATA_SIZE = 64;
								localparam _param_D5D25_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
								if (1) begin : l1_mem_arb_bus_if
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_D5D25_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_D5D25_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:7:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_mem_bus_if.sv:9:5
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:21:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire [612:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire [518:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:30:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:31:5
									// Trace: src/VX_mem_bus_if.sv:39:5
								end
								// Trace: src/VX_socket.sv:232:5
								assign l1_mem_arb_bus_if.req_valid = dcache_mem_bus_if[i].req_valid;
								// Trace: src/VX_socket.sv:233:5
								assign l1_mem_arb_bus_if.req_data[612] = dcache_mem_bus_if[i].req_data[611];
								// Trace: src/VX_socket.sv:234:5
								assign l1_mem_arb_bus_if.req_data[611-:26] = dcache_mem_bus_if[i].req_data[610-:26];
								// Trace: src/VX_socket.sv:235:5
								assign l1_mem_arb_bus_if.req_data[585-:512] = dcache_mem_bus_if[i].req_data[584-:512];
								// Trace: src/VX_socket.sv:236:5
								assign l1_mem_arb_bus_if.req_data[73-:64] = dcache_mem_bus_if[i].req_data[72-:64];
								// Trace: src/VX_socket.sv:237:5
								assign l1_mem_arb_bus_if.req_data[9-:3] = dcache_mem_bus_if[i].req_data[8-:3];
								if (1) begin : genblk1
									if (1) begin : genblk1
										if (1) begin : genblk1
											// Trace: src/VX_socket.sv:242:17
											assign l1_mem_arb_bus_if.req_data[6-:7] = {dcache_mem_bus_if[i].req_data[5-:1], 1'b0, dcache_mem_bus_if[i].req_data[4-:5]};
										end
									end
								end
								// Trace: src/VX_socket.sv:257:5
								assign dcache_mem_bus_if[i].req_ready = l1_mem_arb_bus_if.req_ready;
								// Trace: src/VX_socket.sv:258:5
								assign dcache_mem_bus_if[i].rsp_valid = l1_mem_arb_bus_if.rsp_valid;
								// Trace: src/VX_socket.sv:259:5
								assign dcache_mem_bus_if[i].rsp_data[517-:512] = l1_mem_arb_bus_if.rsp_data[518-:512];
								if (1) begin : genblk2
									if (1) begin : genblk1
										if (1) begin : genblk1
											// Trace: src/VX_socket.sv:264:17
											assign dcache_mem_bus_if[i].rsp_data[5-:6] = {l1_mem_arb_bus_if.rsp_data[6-:1], l1_mem_arb_bus_if.rsp_data[4:0]};
										end
									end
								end
								// Trace: src/VX_socket.sv:279:5
								assign l1_mem_arb_bus_if.rsp_ready = dcache_mem_bus_if[i].rsp_ready;
								// Trace: src/VX_socket.sv:280:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].req_valid = l1_mem_arb_bus_if.req_valid;
								// Trace: src/VX_socket.sv:281:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].req_data = l1_mem_arb_bus_if.req_data;
								// Trace: src/VX_socket.sv:282:5
								assign l1_mem_arb_bus_if.req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
								// Trace: src/VX_socket.sv:283:5
								assign l1_mem_arb_bus_if.rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
								// Trace: src/VX_socket.sv:284:5
								assign l1_mem_arb_bus_if.rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
								// Trace: src/VX_socket.sv:285:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = l1_mem_arb_bus_if.rsp_ready;
							end
						end
						// Trace: src/VX_socket.sv:288:5
						wire [0:0] per_core_busy;
						// Trace: src/VX_socket.sv:289:5
						genvar _gv_core_id_1;
						for (_gv_core_id_1 = 0; _gv_core_id_1 < 1; _gv_core_id_1 = _gv_core_id_1 + 1) begin : g_cores
							localparam core_id = _gv_core_id_1;
							// Trace: src/VX_socket.sv:290:5
							wire [0:0] core_reset;
							// Trace: src/VX_socket.sv:291:5
							VX_reset_relay #(
								.N(1),
								.MAX_FANOUT(0)
							) __core_reset(
								.clk(clk),
								.reset(reset),
								.reset_o(core_reset)
							);
							// Trace: src/VX_socket.sv:296:9
							// expanded interface instance: core_dcr_bus_if
							if (1) begin : core_dcr_bus_if
								// Trace: src/VX_dcr_bus_if.sv:2:5
								wire write_valid;
								// Trace: src/VX_dcr_bus_if.sv:3:5
								wire [11:0] write_addr;
								// Trace: src/VX_dcr_bus_if.sv:4:5
								wire [31:0] write_data;
								// Trace: src/VX_dcr_bus_if.sv:5:5
								// Trace: src/VX_dcr_bus_if.sv:10:5
							end
							if (1) begin : genblk1
								// Trace: src/VX_socket.sv:310:9
								assign {core_dcr_bus_if.write_valid, core_dcr_bus_if.write_addr, core_dcr_bus_if.write_data} = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket_dcr_bus_if.write_valid && 1'b1, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket_dcr_bus_if.write_addr, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket_dcr_bus_if.write_data};
							end
							// Trace: src/VX_socket.sv:313:9
							// expanded module instance: core
							localparam _bbase_588EE_dcache_bus_if = core_id * VX_gpu_pkg_DCACHE_NUM_REQS;
							localparam _bbase_588EE_icache_bus_if = core_id;
							localparam _param_588EE_CORE_ID = (SOCKET_ID * 1) + core_id;
							localparam _param_588EE_INSTANCE_ID = "";
							if (1) begin : core
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_core.sv:2:15
								localparam CORE_ID = _param_588EE_CORE_ID;
								// Trace: src/VX_core.sv:3:16
								localparam INSTANCE_ID = _param_588EE_INSTANCE_ID;
								// Trace: src/VX_core.sv:5:5
								wire clk;
								// Trace: src/VX_core.sv:6:5
								wire reset;
								// Trace: src/VX_core.sv:7:5
								// removed modport instance dcr_bus_if
								// Trace: src/VX_core.sv:8:5
								localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
								localparam VX_gpu_pkg_LSU_WORD_SIZE = 4;
								localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
								localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
								localparam _mbase_dcache_bus_if = _bbase_588EE_dcache_bus_if;
								// Trace: src/VX_core.sv:9:5
								localparam _mbase_icache_bus_if = _bbase_588EE_icache_bus_if;
								// Trace: src/VX_core.sv:10:5
								wire busy;
								// Trace: src/VX_core.sv:12:5
								// expanded interface instance: schedule_if
								if (1) begin : schedule_if
									// Trace: src/VX_schedule_if.sv:2:5
									// removed localparam type data_t
									// Trace: src/VX_schedule_if.sv:8:5
									wire valid;
									// Trace: src/VX_schedule_if.sv:9:5
									wire [37:0] data;
									// Trace: src/VX_schedule_if.sv:10:5
									wire ready;
									// Trace: src/VX_schedule_if.sv:11:5
									// Trace: src/VX_schedule_if.sv:16:5
								end
								// Trace: src/VX_core.sv:13:5
								// expanded interface instance: fetch_if
								if (1) begin : fetch_if
									// Trace: src/VX_fetch_if.sv:2:5
									// removed localparam type data_t
									// Trace: src/VX_fetch_if.sv:9:5
									wire valid;
									// Trace: src/VX_fetch_if.sv:10:5
									wire [69:0] data;
									// Trace: src/VX_fetch_if.sv:11:5
									wire ready;
									// Trace: src/VX_fetch_if.sv:12:5
									// Trace: src/VX_fetch_if.sv:17:5
								end
								// Trace: src/VX_core.sv:14:5
								// expanded interface instance: decode_if
								if (1) begin : decode_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_decode_if.sv:2:15
									localparam NUM_WARPS = 4;
									// Trace: src/VX_decode_if.sv:3:15
									localparam NW_WIDTH = 2;
									// Trace: src/VX_decode_if.sv:5:5
									// removed localparam type VX_gpu_pkg_alu_args_t
									// removed localparam type VX_gpu_pkg_csr_args_t
									// removed localparam type VX_gpu_pkg_fpu_args_t
									// removed localparam type VX_gpu_pkg_lsu_args_t
									// removed localparam type VX_gpu_pkg_wctl_args_t
									// removed localparam type VX_gpu_pkg_op_args_t
									// removed localparam type data_t
									// Trace: src/VX_decode_if.sv:19:5
									wire valid;
									// Trace: src/VX_decode_if.sv:20:5
									wire [105:0] data;
									// Trace: src/VX_decode_if.sv:21:5
									wire ready;
									// Trace: src/VX_decode_if.sv:22:5
									// Trace: src/VX_decode_if.sv:27:5
								end
								// Trace: src/VX_core.sv:15:5
								// expanded interface instance: sched_csr_if
								if (1) begin : sched_csr_if
									// Trace: src/VX_sched_csr_if.sv:2:5
									wire [43:0] cycles;
									// Trace: src/VX_sched_csr_if.sv:3:5
									wire [3:0] active_warps;
									// Trace: src/VX_sched_csr_if.sv:4:5
									wire [15:0] thread_masks;
									// Trace: src/VX_sched_csr_if.sv:5:5
									wire alm_empty;
									// Trace: src/VX_sched_csr_if.sv:6:5
									wire [1:0] alm_empty_wid;
									// Trace: src/VX_sched_csr_if.sv:7:5
									wire unlock_warp;
									// Trace: src/VX_sched_csr_if.sv:8:5
									wire [1:0] unlock_wid;
									// Trace: src/VX_sched_csr_if.sv:9:5
									// Trace: src/VX_sched_csr_if.sv:18:5
								end
								// Trace: src/VX_core.sv:16:5
								// expanded interface instance: decode_sched_if
								if (1) begin : decode_sched_if
									// Trace: src/VX_decode_sched_if.sv:2:5
									wire valid;
									// Trace: src/VX_decode_sched_if.sv:3:5
									wire unlock;
									// Trace: src/VX_decode_sched_if.sv:4:5
									wire [1:0] wid;
									// Trace: src/VX_decode_sched_if.sv:5:5
									// Trace: src/VX_decode_sched_if.sv:10:5
								end
								// Trace: src/VX_core.sv:17:5
								// expanded interface instance: commit_sched_if
								if (1) begin : commit_sched_if
									// Trace: src/VX_commit_sched_if.sv:2:5
									wire [3:0] committed_warps;
									// Trace: src/VX_commit_sched_if.sv:3:5
									// Trace: src/VX_commit_sched_if.sv:6:5
								end
								// Trace: src/VX_core.sv:18:5
								// expanded interface instance: commit_csr_if
								if (1) begin : commit_csr_if
									// Trace: src/VX_commit_csr_if.sv:2:5
									wire [43:0] instret;
									// Trace: src/VX_commit_csr_if.sv:3:5
									// Trace: src/VX_commit_csr_if.sv:6:5
								end
								// Trace: src/VX_core.sv:19:5
								// expanded interface instance: branch_ctl_if
								genvar _arr_DDFE6;
								for (_arr_DDFE6 = 0; _arr_DDFE6 <= 0; _arr_DDFE6 = _arr_DDFE6 + 1) begin : branch_ctl_if
									// Trace: src/VX_branch_ctl_if.sv:2:5
									wire valid;
									// Trace: src/VX_branch_ctl_if.sv:3:5
									wire [1:0] wid;
									// Trace: src/VX_branch_ctl_if.sv:4:5
									wire taken;
									// Trace: src/VX_branch_ctl_if.sv:5:5
									wire [30:0] dest;
									// Trace: src/VX_branch_ctl_if.sv:6:5
									// Trace: src/VX_branch_ctl_if.sv:12:5
								end
								// Trace: src/VX_core.sv:20:5
								// expanded interface instance: warp_ctl_if
								if (1) begin : warp_ctl_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_warp_ctl_if.sv:2:5
									wire valid;
									// Trace: src/VX_warp_ctl_if.sv:3:5
									wire [1:0] wid;
									// Trace: src/VX_warp_ctl_if.sv:4:5
									// removed localparam type VX_gpu_pkg_tmc_t
									wire [4:0] tmc;
									// Trace: src/VX_warp_ctl_if.sv:5:5
									// removed localparam type VX_gpu_pkg_wspawn_t
									wire [35:0] wspawn;
									// Trace: src/VX_warp_ctl_if.sv:6:5
									// removed localparam type VX_gpu_pkg_split_t
									wire [40:0] split;
									// Trace: src/VX_warp_ctl_if.sv:7:5
									// removed localparam type VX_gpu_pkg_join_t
									wire [2:0] sjoin;
									// Trace: src/VX_warp_ctl_if.sv:8:5
									// removed localparam type VX_gpu_pkg_barrier_t
									wire [5:0] barrier;
									// Trace: src/VX_warp_ctl_if.sv:9:5
									wire [1:0] dvstack_wid;
									// Trace: src/VX_warp_ctl_if.sv:10:5
									wire [1:0] dvstack_ptr;
									// Trace: src/VX_warp_ctl_if.sv:11:5
									// Trace: src/VX_warp_ctl_if.sv:22:5
								end
								// Trace: src/VX_core.sv:21:5
								// expanded interface instance: dispatch_if
								genvar _arr_B1D72;
								for (_arr_B1D72 = 0; _arr_B1D72 <= 3; _arr_B1D72 = _arr_B1D72 + 1) begin : dispatch_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_dispatch_if.sv:2:5
									localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
									localparam VX_gpu_pkg_ISSUE_WIS = 2;
									localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
									// removed localparam type VX_gpu_pkg_alu_args_t
									// removed localparam type VX_gpu_pkg_csr_args_t
									// removed localparam type VX_gpu_pkg_fpu_args_t
									// removed localparam type VX_gpu_pkg_lsu_args_t
									// removed localparam type VX_gpu_pkg_wctl_args_t
									// removed localparam type VX_gpu_pkg_op_args_t
									// removed localparam type data_t
									// Trace: src/VX_dispatch_if.sv:16:5
									wire valid;
									// Trace: src/VX_dispatch_if.sv:17:5
									wire [471:0] data;
									// Trace: src/VX_dispatch_if.sv:18:5
									wire ready;
									// Trace: src/VX_dispatch_if.sv:19:5
									// Trace: src/VX_dispatch_if.sv:24:5
								end
								// Trace: src/VX_core.sv:22:5
								// expanded interface instance: commit_if
								genvar _arr_56FA2;
								for (_arr_56FA2 = 0; _arr_56FA2 <= 3; _arr_56FA2 = _arr_56FA2 + 1) begin : commit_if
									// Trace: src/VX_commit_if.sv:2:15
									localparam NUM_LANES = 4;
									// Trace: src/VX_commit_if.sv:3:15
									localparam PID_WIDTH = 1;
									// Trace: src/VX_commit_if.sv:5:5
									// removed localparam type data_t
									// Trace: src/VX_commit_if.sv:17:5
									wire valid;
									// Trace: src/VX_commit_if.sv:18:5
									wire [175:0] data;
									// Trace: src/VX_commit_if.sv:19:5
									wire ready;
									// Trace: src/VX_commit_if.sv:20:5
									// Trace: src/VX_commit_if.sv:25:5
								end
								// Trace: src/VX_core.sv:23:5
								// expanded interface instance: writeback_if
								genvar _arr_8BCF0;
								for (_arr_8BCF0 = 0; _arr_8BCF0 <= 0; _arr_8BCF0 = _arr_8BCF0 + 1) begin : writeback_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_writeback_if.sv:2:5
									localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
									localparam VX_gpu_pkg_ISSUE_WIS = 2;
									localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
									// removed localparam type data_t
									// Trace: src/VX_writeback_if.sv:12:5
									wire valid;
									// Trace: src/VX_writeback_if.sv:13:5
									wire [173:0] data;
									// Trace: src/VX_writeback_if.sv:14:5
									// Trace: src/VX_writeback_if.sv:18:5
								end
								// Trace: src/VX_core.sv:24:5
								localparam VX_gpu_pkg_LSU_MEM_BATCHES = 1;
								localparam VX_gpu_pkg_LSU_TAG_ID_BITS = 1;
								localparam VX_gpu_pkg_LSU_TAG_WIDTH = 2;
								// expanded interface instance: lsu_mem_if
								localparam _param_DD8FC_NUM_LANES = 4;
								localparam _param_DD8FC_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
								localparam _param_DD8FC_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
								genvar _arr_DD8FC;
								for (_arr_DD8FC = 0; _arr_DD8FC <= 0; _arr_DD8FC = _arr_DD8FC + 1) begin : lsu_mem_if
									// Trace: src/VX_lsu_mem_if.sv:2:15
									localparam NUM_LANES = _param_DD8FC_NUM_LANES;
									// Trace: src/VX_lsu_mem_if.sv:3:15
									localparam DATA_SIZE = _param_DD8FC_DATA_SIZE;
									// Trace: src/VX_lsu_mem_if.sv:4:15
									localparam TAG_WIDTH = _param_DD8FC_TAG_WIDTH;
									// Trace: src/VX_lsu_mem_if.sv:5:15
									localparam FLAGS_WIDTH = 3;
									// Trace: src/VX_lsu_mem_if.sv:6:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_lsu_mem_if.sv:7:15
									localparam ADDR_WIDTH = 30;
									// Trace: src/VX_lsu_mem_if.sv:8:15
									localparam UUID_WIDTH = 1;
									// Trace: src/VX_lsu_mem_if.sv:10:5
									// removed localparam type tag_t
									// Trace: src/VX_lsu_mem_if.sv:14:5
									// removed localparam type req_data_t
									// Trace: src/VX_lsu_mem_if.sv:23:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_lsu_mem_if.sv:28:5
									wire req_valid;
									// Trace: src/VX_lsu_mem_if.sv:29:5
									wire [282:0] req_data;
									// Trace: src/VX_lsu_mem_if.sv:30:5
									wire req_ready;
									// Trace: src/VX_lsu_mem_if.sv:31:5
									wire rsp_valid;
									// Trace: src/VX_lsu_mem_if.sv:32:5
									wire [133:0] rsp_data;
									// Trace: src/VX_lsu_mem_if.sv:33:5
									wire rsp_ready;
									// Trace: src/VX_lsu_mem_if.sv:34:5
									// Trace: src/VX_lsu_mem_if.sv:42:5
								end
								// Trace: src/VX_core.sv:29:5
								// removed localparam type VX_gpu_pkg_base_dcrs_t
								wire [71:0] base_dcrs;
								// Trace: src/VX_core.sv:30:5
								// expanded module instance: dcr_data
								if (1) begin : dcr_data
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_dcr_data.sv:2:5
									wire clk;
									// Trace: src/VX_dcr_data.sv:3:5
									wire reset;
									// Trace: src/VX_dcr_data.sv:4:5
									// removed modport instance dcr_bus_if
									// Trace: src/VX_dcr_data.sv:5:5
									// removed localparam type VX_gpu_pkg_base_dcrs_t
									wire [71:0] base_dcrs;
									// Trace: src/VX_dcr_data.sv:7:5
									reg [71:0] dcrs;
									// Trace: src/VX_dcr_data.sv:8:5
									always @(posedge clk)
										// Trace: src/VX_dcr_data.sv:9:8
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_valid)
											// Trace: src/VX_dcr_data.sv:10:13
											case (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_addr)
												12'h001:
													// Trace: src/VX_dcr_data.sv:11:23
													dcrs[71:40] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_data;
												12'h003:
													// Trace: src/VX_dcr_data.sv:12:23
													dcrs[39:8] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_data;
												12'h005:
													// Trace: src/VX_dcr_data.sv:13:23
													dcrs[7-:8] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_data[7:0];
												default:
													;
											endcase
									// Trace: src/VX_dcr_data.sv:18:5
									assign base_dcrs = dcrs;
								end
								assign dcr_data.clk = clk;
								assign dcr_data.reset = reset;
								assign base_dcrs = dcr_data.base_dcrs;
								// Trace: src/VX_core.sv:37:5
								// expanded module instance: schedule
								localparam _bbase_45092_branch_ctl_if = 0;
								localparam _param_45092_INSTANCE_ID = "";
								localparam _param_45092_CORE_ID = CORE_ID;
								if (1) begin : schedule
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_schedule.sv:2:16
									localparam INSTANCE_ID = _param_45092_INSTANCE_ID;
									// Trace: src/VX_schedule.sv:3:15
									localparam CORE_ID = _param_45092_CORE_ID;
									// Trace: src/VX_schedule.sv:5:5
									wire clk;
									// Trace: src/VX_schedule.sv:6:5
									wire reset;
									// Trace: src/VX_schedule.sv:7:5
									// removed localparam type VX_gpu_pkg_base_dcrs_t
									wire [71:0] base_dcrs;
									// Trace: src/VX_schedule.sv:8:5
									// removed modport instance warp_ctl_if
									// Trace: src/VX_schedule.sv:9:5
									localparam _mbase_branch_ctl_if = 0;
									// Trace: src/VX_schedule.sv:10:5
									// removed modport instance decode_sched_if
									// Trace: src/VX_schedule.sv:11:5
									// removed modport instance commit_sched_if
									// Trace: src/VX_schedule.sv:12:5
									// removed modport instance schedule_if
									// Trace: src/VX_schedule.sv:13:5
									// removed modport instance sched_csr_if
									// Trace: src/VX_schedule.sv:14:5
									wire busy;
									// Trace: src/VX_schedule.sv:16:5
									reg [3:0] active_warps;
									reg [3:0] active_warps_n;
									// Trace: src/VX_schedule.sv:17:5
									reg [3:0] stalled_warps;
									reg [3:0] stalled_warps_n;
									// Trace: src/VX_schedule.sv:18:5
									reg [15:0] thread_masks;
									reg [15:0] thread_masks_n;
									// Trace: src/VX_schedule.sv:19:5
									reg [123:0] warp_pcs;
									reg [123:0] warp_pcs_n;
									// Trace: src/VX_schedule.sv:20:5
									wire [1:0] schedule_wid;
									// Trace: src/VX_schedule.sv:21:5
									wire [3:0] schedule_tmask;
									// Trace: src/VX_schedule.sv:22:5
									wire [30:0] schedule_pc;
									// Trace: src/VX_schedule.sv:23:5
									wire schedule_valid;
									// Trace: src/VX_schedule.sv:24:5
									wire schedule_ready;
									// Trace: src/VX_schedule.sv:25:5
									wire join_valid;
									// Trace: src/VX_schedule.sv:26:5
									wire join_is_dvg;
									// Trace: src/VX_schedule.sv:27:5
									wire join_is_else;
									// Trace: src/VX_schedule.sv:28:5
									wire [1:0] join_wid;
									// Trace: src/VX_schedule.sv:29:5
									wire [3:0] join_tmask;
									// Trace: src/VX_schedule.sv:30:5
									wire [30:0] join_pc;
									// Trace: src/VX_schedule.sv:31:5
									reg [43:0] cycles;
									// Trace: src/VX_schedule.sv:32:5
									reg [3:0] issued_instrs;
									// Trace: src/VX_schedule.sv:33:5
									wire schedule_fire = schedule_valid && schedule_ready;
									// Trace: src/VX_schedule.sv:34:5
									wire schedule_if_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.ready;
									// Trace: src/VX_schedule.sv:35:5
									wire [0:0] branch_valid;
									// Trace: src/VX_schedule.sv:36:5
									wire [1:0] branch_wid;
									// Trace: src/VX_schedule.sv:37:5
									wire [0:0] branch_taken;
									// Trace: src/VX_schedule.sv:38:5
									wire [30:0] branch_dest;
									// Trace: src/VX_schedule.sv:39:5
									genvar _gv_i_145;
									for (_gv_i_145 = 0; _gv_i_145 < 1; _gv_i_145 = _gv_i_145 + 1) begin : g_branch_init
										localparam i = _gv_i_145;
										// Trace: src/VX_schedule.sv:40:9
										assign branch_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[i + _mbase_branch_ctl_if].valid;
										// Trace: src/VX_schedule.sv:41:9
										assign branch_wid[i * 2+:2] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[i + _mbase_branch_ctl_if].wid;
										// Trace: src/VX_schedule.sv:42:9
										assign branch_taken[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[i + _mbase_branch_ctl_if].taken;
										// Trace: src/VX_schedule.sv:43:9
										assign branch_dest[i * 31+:31] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[i + _mbase_branch_ctl_if].dest;
									end
									// Trace: src/VX_schedule.sv:45:5
									reg [7:0] barrier_masks;
									reg [7:0] barrier_masks_n;
									// Trace: src/VX_schedule.sv:46:5
									reg [3:0] barrier_ctrs;
									reg [3:0] barrier_ctrs_n;
									// Trace: src/VX_schedule.sv:47:5
									reg [3:0] barrier_stalls;
									reg [3:0] barrier_stalls_n;
									// Trace: src/VX_schedule.sv:48:5
									reg [3:0] curr_barrier_mask_p1;
									// Trace: src/VX_schedule.sv:49:5
									// removed localparam type VX_gpu_pkg_wspawn_t
									reg [35:0] wspawn;
									// Trace: src/VX_schedule.sv:50:5
									reg [1:0] wspawn_wid;
									// Trace: src/VX_schedule.sv:51:5
									reg is_single_warp;
									// Trace: src/VX_schedule.sv:52:5
									wire [2:0] active_warps_cnt;
									// Trace: src/VX_schedule.sv:53:5
									VX_popcount #(
										.N(4),
										.MODEL(1)
									) __active_warps_cnt__(
										.data_in(active_warps),
										.data_out(active_warps_cnt)
									);
									// Trace: src/VX_schedule.sv:60:5
									always @(*) begin
										// Trace: src/VX_schedule.sv:61:9
										active_warps_n = active_warps;
										// Trace: src/VX_schedule.sv:62:9
										stalled_warps_n = stalled_warps;
										// Trace: src/VX_schedule.sv:63:9
										thread_masks_n = thread_masks;
										// Trace: src/VX_schedule.sv:64:9
										barrier_masks_n = barrier_masks;
										// Trace: src/VX_schedule.sv:65:9
										barrier_ctrs_n = barrier_ctrs;
										// Trace: src/VX_schedule.sv:66:9
										barrier_stalls_n = barrier_stalls;
										// Trace: src/VX_schedule.sv:67:9
										warp_pcs_n = warp_pcs;
										// Trace: src/VX_schedule.sv:68:9
										if (wspawn[35] && is_single_warp) begin
											// Trace: src/VX_schedule.sv:69:13
											active_warps_n = active_warps_n | wspawn[34-:4];
											// Trace: src/VX_schedule.sv:70:13
											begin : sv2v_autoblock_3
												// Trace: src/VX_schedule.sv:70:18
												integer i;
												// Trace: src/VX_schedule.sv:70:18
												for (i = 0; i < 4; i = i + 1)
													begin
														// Trace: src/VX_schedule.sv:71:17
														if (wspawn[31 + i]) begin
															// Trace: src/VX_schedule.sv:72:21
															thread_masks_n[i * 4] = 1;
															// Trace: src/VX_schedule.sv:73:21
															warp_pcs_n[i * 31+:31] = wspawn[30-:31];
														end
													end
											end
											// Trace: src/VX_schedule.sv:76:13
											stalled_warps_n[wspawn_wid] = 0;
										end
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.tmc[4]) begin
											// Trace: src/VX_schedule.sv:79:13
											active_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.tmc[3-:4] != 0;
											// Trace: src/VX_schedule.sv:80:13
											thread_masks_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid * 4+:4] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.tmc[3-:4];
											// Trace: src/VX_schedule.sv:81:13
											stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 0;
										end
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split[40]) begin
											// Trace: src/VX_schedule.sv:84:13
											if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split[39])
												// Trace: src/VX_schedule.sv:85:17
												thread_masks_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid * 4+:4] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split[38-:4];
											// Trace: src/VX_schedule.sv:87:13
											stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 0;
										end
										if (join_valid) begin
											// Trace: src/VX_schedule.sv:90:13
											if (join_is_dvg) begin
												// Trace: src/VX_schedule.sv:91:17
												if (join_is_else)
													// Trace: src/VX_schedule.sv:92:21
													warp_pcs_n[join_wid * 31+:31] = join_pc;
												// Trace: src/VX_schedule.sv:94:17
												thread_masks_n[join_wid * 4+:4] = join_tmask;
											end
											// Trace: src/VX_schedule.sv:96:13
											stalled_warps_n[join_wid] = 0;
										end
										// Trace: src/VX_schedule.sv:98:9
										curr_barrier_mask_p1 = barrier_masks[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 4+:4];
										// Trace: src/VX_schedule.sv:99:9
										curr_barrier_mask_p1[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 1;
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[5]) begin
											begin
												// Trace: src/VX_schedule.sv:101:13
												if (~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[0]) begin
													begin
														// Trace: src/VX_schedule.sv:102:17
														if (~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[3] && (barrier_ctrs[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 2+:2] == sv2v_cast_2(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[2-:2]))) begin
															// Trace: src/VX_schedule.sv:104:21
															barrier_ctrs_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 2+:2] = 1'sb0;
															// Trace: src/VX_schedule.sv:105:21
															barrier_masks_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 4+:4] = 1'sb0;
															// Trace: src/VX_schedule.sv:106:21
															stalled_warps_n = stalled_warps_n & ~barrier_masks[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 4+:4];
															// Trace: src/VX_schedule.sv:107:21
															stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 0;
														end
														else begin
															// Trace: src/VX_schedule.sv:109:21
															barrier_ctrs_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 2+:2] = barrier_ctrs[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 2+:2] + 2'sd1;
															// Trace: src/VX_schedule.sv:110:21
															barrier_masks_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 4+:4] = curr_barrier_mask_p1;
														end
													end
												end
												else
													// Trace: src/VX_schedule.sv:113:17
													stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 0;
											end
										end
										begin : sv2v_autoblock_4
											// Trace: src/VX_schedule.sv:116:14
											integer i;
											// Trace: src/VX_schedule.sv:116:14
											for (i = 0; i < 1; i = i + 1)
												begin
													// Trace: src/VX_schedule.sv:117:13
													if (branch_valid[i]) begin
														// Trace: src/VX_schedule.sv:118:17
														if (branch_taken[i])
															// Trace: src/VX_schedule.sv:119:21
															warp_pcs_n[branch_wid[i * 2+:2] * 31+:31] = branch_dest[i * 31+:31];
														// Trace: src/VX_schedule.sv:121:17
														stalled_warps_n[branch_wid[i * 2+:2]] = 0;
													end
												end
										end
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.unlock)
											// Trace: src/VX_schedule.sv:125:13
											stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.wid] = 0;
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.unlock_warp)
											// Trace: src/VX_schedule.sv:128:13
											stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.unlock_wid] = 0;
										if (schedule_fire)
											// Trace: src/VX_schedule.sv:131:13
											stalled_warps_n[schedule_wid] = 1;
										if (schedule_if_fire)
											// Trace: src/VX_schedule.sv:134:13
											warp_pcs_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[36-:2] * 31+:31] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[30-:31] + 31'sd2;
									end
									// Trace: src/VX_schedule.sv:137:5
									always @(posedge clk)
										// Trace: src/VX_schedule.sv:138:9
										if (reset) begin
											// Trace: src/VX_schedule.sv:139:13
											barrier_masks <= 1'sb0;
											// Trace: src/VX_schedule.sv:140:13
											barrier_ctrs <= 1'sb0;
											// Trace: src/VX_schedule.sv:141:13
											stalled_warps <= 1'sb0;
											// Trace: src/VX_schedule.sv:142:13
											warp_pcs <= 1'sb0;
											// Trace: src/VX_schedule.sv:143:13
											active_warps <= 1'sb0;
											// Trace: src/VX_schedule.sv:144:13
											thread_masks <= 1'sb0;
											// Trace: src/VX_schedule.sv:145:13
											barrier_stalls <= 1'sb0;
											// Trace: src/VX_schedule.sv:146:13
											issued_instrs <= 1'sb0;
											// Trace: src/VX_schedule.sv:147:13
											cycles <= 1'sb0;
											// Trace: src/VX_schedule.sv:148:13
											wspawn[35] <= 0;
											// Trace: src/VX_schedule.sv:149:13
											warp_pcs[0+:31] <= base_dcrs[41+:31];
											// Trace: src/VX_schedule.sv:150:13
											active_warps[0] <= 1;
											// Trace: src/VX_schedule.sv:151:13
											thread_masks[0] <= 1;
											// Trace: src/VX_schedule.sv:152:13
											is_single_warp <= 1;
										end
										else begin
											// Trace: src/VX_schedule.sv:154:13
											active_warps <= active_warps_n;
											// Trace: src/VX_schedule.sv:155:13
											stalled_warps <= stalled_warps_n;
											// Trace: src/VX_schedule.sv:156:13
											thread_masks <= thread_masks_n;
											// Trace: src/VX_schedule.sv:157:13
											warp_pcs <= warp_pcs_n;
											// Trace: src/VX_schedule.sv:158:13
											barrier_masks <= barrier_masks_n;
											// Trace: src/VX_schedule.sv:159:13
											barrier_ctrs <= barrier_ctrs_n;
											// Trace: src/VX_schedule.sv:160:13
											barrier_stalls <= barrier_stalls_n;
											// Trace: src/VX_schedule.sv:161:13
											is_single_warp <= active_warps_cnt == sv2v_cast_22555_signed(1);
											// Trace: src/VX_schedule.sv:162:13
											if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wspawn[35]) begin
												// Trace: src/VX_schedule.sv:163:17
												wspawn[35] <= 1;
												// Trace: src/VX_schedule.sv:164:17
												wspawn[34-:4] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wspawn[34-:4];
												// Trace: src/VX_schedule.sv:165:17
												wspawn[30-:31] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wspawn[30-:31];
												// Trace: src/VX_schedule.sv:166:17
												wspawn_wid <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid;
											end
											if (wspawn[35] && is_single_warp)
												// Trace: src/VX_schedule.sv:169:17
												wspawn[35] <= 0;
											if (schedule_if_fire)
												// Trace: src/VX_schedule.sv:172:17
												issued_instrs[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[36-:2]+:1] <= issued_instrs[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[36-:2]+:1] + 1'sd1;
											if (busy)
												// Trace: src/VX_schedule.sv:175:17
												cycles <= cycles + 1;
										end
									// Trace: src/VX_schedule.sv:179:5
									VX_split_join #(.INSTANCE_ID("")) split_join(
										.clk(clk),
										.reset(reset),
										.valid(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid),
										.wid(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid),
										.split(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split),
										.sjoin(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.sjoin),
										.join_valid(join_valid),
										.join_is_dvg(join_is_dvg),
										.join_is_else(join_is_else),
										.join_wid(join_wid),
										.join_tmask(join_tmask),
										.join_pc(join_pc),
										.stack_wid(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.dvstack_wid),
										.stack_ptr(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.dvstack_ptr)
									);
									// Trace: src/VX_schedule.sv:197:5
									wire [3:0] ready_warps = active_warps & ~stalled_warps;
									// Trace: src/VX_schedule.sv:198:5
									VX_lzc #(
										.N(4),
										.REVERSE(1)
									) wid_select(
										.data_in(ready_warps),
										.data_out(schedule_wid),
										.valid_out(schedule_valid)
									);
									// Trace: src/VX_schedule.sv:206:5
									wire [139:0] schedule_data;
									// Trace: src/VX_schedule.sv:207:5
									genvar _gv_i_146;
									for (_gv_i_146 = 0; _gv_i_146 < 4; _gv_i_146 = _gv_i_146 + 1) begin : g_schedule_data
										localparam i = _gv_i_146;
										// Trace: src/VX_schedule.sv:208:9
										assign schedule_data[i * 35+:35] = {thread_masks[i * 4+:4], warp_pcs[i * 31+:31]};
									end
									// Trace: src/VX_schedule.sv:210:5
									assign {schedule_tmask, schedule_pc} = {schedule_data[(schedule_wid * 35) + 34-:4], schedule_data[(schedule_wid * 35) + 30-:31]};
									// Trace: src/VX_schedule.sv:214:5
									wire [0:0] instr_uuid;
									// Trace: src/VX_schedule.sv:215:5
									assign instr_uuid = 1'sb0;
									// Trace: src/VX_schedule.sv:216:5
									VX_elastic_buffer #(
										.DATAW(38),
										.SIZE(2),
										.OUT_REG(1)
									) out_buf(
										.clk(clk),
										.reset(reset),
										.valid_in(schedule_valid),
										.ready_in(schedule_ready),
										.data_in({schedule_tmask, schedule_pc, schedule_wid, instr_uuid}),
										.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[34-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[30-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[36-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[37]}),
										.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.valid),
										.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.ready)
									);
									// Trace: src/VX_schedule.sv:230:5
									wire [3:0] pending_warp_empty;
									// Trace: src/VX_schedule.sv:231:5
									wire [3:0] pending_warp_alm_empty;
									// Trace: src/VX_schedule.sv:232:5
									genvar _gv_i_147;
									for (_gv_i_147 = 0; _gv_i_147 < 4; _gv_i_147 = _gv_i_147 + 1) begin : g_pending_sizes
										localparam i = _gv_i_147;
										// Trace: src/VX_schedule.sv:233:9
										VX_pending_size #(
											.SIZE(4096),
											.ALM_EMPTY(1)
										) counter(
											.clk(clk),
											.reset(reset),
											.incr(schedule_if_fire && (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[36-:2] == sv2v_cast_2_signed(i))),
											.decr(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_sched_if.committed_warps[i]),
											.empty(pending_warp_empty[i]),
											.alm_empty(pending_warp_alm_empty[i]),
											.full(),
											.alm_full(),
											.size()
										);
									end
									// Trace: src/VX_schedule.sv:248:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.alm_empty = pending_warp_alm_empty[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.alm_empty_wid];
									// Trace: src/VX_schedule.sv:249:5
									wire no_pending_instr = &pending_warp_empty;
									// Trace: src/VX_schedule.sv:250:5
									VX_pipe_register #(
										.DATAW(1),
										.RESETW(1),
										.DEPTH(1)
									) __busy__(
										.clk(clk),
										.reset(reset),
										.enable(1'b1),
										.data_in((active_warps != 0) || ~no_pending_instr),
										.data_out(busy)
									);
									// Trace: src/VX_schedule.sv:261:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.cycles = cycles;
									// Trace: src/VX_schedule.sv:262:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.active_warps = active_warps;
									// Trace: src/VX_schedule.sv:263:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.thread_masks = thread_masks;
									// Trace: src/VX_schedule.sv:264:5
									reg [31:0] timeout_ctr;
									// Trace: src/VX_schedule.sv:265:5
									reg timeout_enable;
									// Trace: src/VX_schedule.sv:266:5
									always @(posedge clk)
										// Trace: src/VX_schedule.sv:267:9
										if (reset) begin
											// Trace: src/VX_schedule.sv:268:13
											timeout_ctr <= 1'sb0;
											// Trace: src/VX_schedule.sv:269:13
											timeout_enable <= 0;
										end
										else begin
											// Trace: src/VX_schedule.sv:271:13
											if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.unlock)
												// Trace: src/VX_schedule.sv:272:17
												timeout_enable <= 1;
											if ((timeout_enable && (active_warps != 0)) && (active_warps == stalled_warps))
												// Trace: src/VX_schedule.sv:275:17
												timeout_ctr <= timeout_ctr + 1;
											else if ((active_warps == 0) || (active_warps != stalled_warps))
												// Trace: src/VX_schedule.sv:277:17
												timeout_ctr <= 1'sb0;
										end
								end
								assign schedule.clk = clk;
								assign schedule.reset = reset;
								assign schedule.base_dcrs = base_dcrs;
								assign busy = schedule.busy;
								// Trace: src/VX_core.sv:52:5
								// expanded module instance: fetch
								localparam _bbase_852F6_icache_bus_if = core_id;
								localparam _param_852F6_INSTANCE_ID = "";
								if (1) begin : fetch
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_fetch.sv:2:16
									localparam INSTANCE_ID = _param_852F6_INSTANCE_ID;
									// Trace: src/VX_fetch.sv:4:5
									wire clk;
									// Trace: src/VX_fetch.sv:5:5
									wire reset;
									// Trace: src/VX_fetch.sv:6:5
									localparam _mbase_icache_bus_if = _bbase_852F6_icache_bus_if;
									// Trace: src/VX_fetch.sv:7:5
									// removed modport instance schedule_if
									// Trace: src/VX_fetch.sv:8:5
									// removed modport instance fetch_if
									// Trace: src/VX_fetch.sv:10:5
									wire icache_req_valid;
									// Trace: src/VX_fetch.sv:11:5
									localparam VX_gpu_pkg_ICACHE_WORD_SIZE = 4;
									localparam VX_gpu_pkg_ICACHE_ADDR_WIDTH = 30;
									wire [29:0] icache_req_addr;
									// Trace: src/VX_fetch.sv:12:5
									localparam VX_gpu_pkg_ICACHE_TAG_ID_BITS = 2;
									localparam VX_gpu_pkg_ICACHE_TAG_WIDTH = 3;
									wire [2:0] icache_req_tag;
									// Trace: src/VX_fetch.sv:13:5
									wire icache_req_ready;
									// Trace: src/VX_fetch.sv:14:5
									wire [0:0] rsp_uuid;
									// Trace: src/VX_fetch.sv:15:5
									wire [1:0] req_tag;
									wire [1:0] rsp_tag;
									// Trace: src/VX_fetch.sv:16:5
									wire icache_req_fire = icache_req_valid && icache_req_ready;
									// Trace: src/VX_fetch.sv:17:5
									assign req_tag = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[36-:2];
									// Trace: src/VX_fetch.sv:18:5
									assign {rsp_uuid, rsp_tag} = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].rsp_data[2-:3];
									// Trace: src/VX_fetch.sv:19:5
									wire [30:0] rsp_PC;
									// Trace: src/VX_fetch.sv:20:5
									wire [3:0] rsp_tmask;
									// Trace: src/VX_fetch.sv:21:5
									VX_dp_ram #(
										.DATAW(35),
										.SIZE(4),
										.RDW_MODE("R")
									) tag_store(
										.clk(clk),
										.reset(reset),
										.read(1'b1),
										.write(icache_req_fire),
										.wren(1'b1),
										.waddr(req_tag),
										.wdata({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[30-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[34-:4]}),
										.raddr(rsp_tag),
										.rdata({rsp_PC, rsp_tmask})
									);
									// Trace: src/VX_fetch.sv:36:5
									wire ibuf_ready = 1'b1;
									// Trace: src/VX_fetch.sv:37:5
									assign icache_req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.valid && ibuf_ready;
									// Trace: src/VX_fetch.sv:38:5
									assign icache_req_addr = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[1+:VX_gpu_pkg_ICACHE_ADDR_WIDTH];
									// Trace: src/VX_fetch.sv:39:5
									assign icache_req_tag = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[37], req_tag};
									// Trace: src/VX_fetch.sv:40:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.ready = icache_req_ready && ibuf_ready;
									// Trace: src/VX_fetch.sv:41:5
									VX_elastic_buffer #(
										.DATAW(33),
										.SIZE(2),
										.OUT_REG(1)
									) req_buf(
										.clk(clk),
										.reset(reset),
										.valid_in(icache_req_valid),
										.ready_in(icache_req_ready),
										.data_in({icache_req_addr, icache_req_tag}),
										.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[71-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[2-:3]}),
										.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_valid),
										.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_ready)
									);
									// Trace: src/VX_fetch.sv:55:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[5-:3] = 1'sb0;
									// Trace: src/VX_fetch.sv:56:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[72] = 0;
									// Trace: src/VX_fetch.sv:57:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[9-:4] = 1'sb1;
									// Trace: src/VX_fetch.sv:58:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[41-:32] = 1'sb0;
									// Trace: src/VX_fetch.sv:59:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].rsp_valid;
									// Trace: src/VX_fetch.sv:60:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[66-:4] = rsp_tmask;
									// Trace: src/VX_fetch.sv:61:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[68-:2] = rsp_tag;
									// Trace: src/VX_fetch.sv:62:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[62-:31] = rsp_PC;
									// Trace: src/VX_fetch.sv:63:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[31-:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].rsp_data[34-:32];
									// Trace: src/VX_fetch.sv:64:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[69] = rsp_uuid;
									// Trace: src/VX_fetch.sv:65:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.ready;
								end
								assign fetch.clk = clk;
								assign fetch.reset = reset;
								// Trace: src/VX_core.sv:61:5
								// expanded module instance: decode
								localparam _param_21B54_INSTANCE_ID = "";
								if (1) begin : decode
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_decode.sv:2:16
									localparam INSTANCE_ID = _param_21B54_INSTANCE_ID;
									// Trace: src/VX_decode.sv:4:5
									wire clk;
									// Trace: src/VX_decode.sv:5:5
									wire reset;
									// Trace: src/VX_decode.sv:6:5
									// removed modport instance fetch_if
									// Trace: src/VX_decode.sv:7:5
									// removed modport instance decode_if
									// Trace: src/VX_decode.sv:8:5
									// removed modport instance decode_sched_if
									// Trace: src/VX_decode.sv:10:5
									// removed localparam type VX_gpu_pkg_alu_args_t
									// removed localparam type VX_gpu_pkg_csr_args_t
									// removed localparam type VX_gpu_pkg_fpu_args_t
									// removed localparam type VX_gpu_pkg_lsu_args_t
									// removed localparam type VX_gpu_pkg_wctl_args_t
									// removed localparam type VX_gpu_pkg_op_args_t
									localparam DATAW = 106;
									// Trace: src/VX_decode.sv:11:5
									reg [1:0] ex_type;
									// Trace: src/VX_decode.sv:12:5
									reg [3:0] op_type;
									// Trace: src/VX_decode.sv:13:5
									reg [36:0] op_args;
									// Trace: src/VX_decode.sv:14:5
									reg [5:0] rd_v;
									reg [5:0] rs1_v;
									reg [5:0] rs2_v;
									reg [5:0] rs3_v;
									// Trace: src/VX_decode.sv:15:5
									reg use_rd;
									reg use_rs1;
									reg use_rs2;
									reg use_rs3;
									// Trace: src/VX_decode.sv:16:5
									reg is_wstall;
									// Trace: src/VX_decode.sv:17:5
									wire [31:0] instr = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[31-:32];
									// Trace: src/VX_decode.sv:18:5
									wire [6:0] opcode = instr[6:0];
									// Trace: src/VX_decode.sv:19:5
									wire [1:0] func2 = instr[26:25];
									// Trace: src/VX_decode.sv:20:5
									wire [2:0] func3 = instr[14:12];
									// Trace: src/VX_decode.sv:21:5
									wire [4:0] func5 = instr[31:27];
									// Trace: src/VX_decode.sv:22:5
									wire [6:0] func7 = instr[31:25];
									// Trace: src/VX_decode.sv:23:5
									wire [11:0] u_12 = instr[31:20];
									// Trace: src/VX_decode.sv:24:5
									wire [4:0] rd = instr[11:7];
									// Trace: src/VX_decode.sv:25:5
									wire [4:0] rs1 = instr[19:15];
									// Trace: src/VX_decode.sv:26:5
									wire [4:0] rs2 = instr[24:20];
									// Trace: src/VX_decode.sv:27:5
									wire [4:0] rs3 = instr[31:27];
									// Trace: src/VX_decode.sv:28:5
									wire is_itype_sh = func3[0] && ~func3[1];
									// Trace: src/VX_decode.sv:29:5
									wire is_fpu_csr = u_12 <= 12'h003;
									// Trace: src/VX_decode.sv:30:5
									wire [19:0] ui_imm = instr[31:12];
									// Trace: src/VX_decode.sv:31:5
									wire [11:0] i_imm = (is_itype_sh ? {7'b0000000, instr[24:20]} : u_12);
									// Trace: src/VX_decode.sv:32:5
									wire [11:0] s_imm = {func7, rd};
									// Trace: src/VX_decode.sv:33:5
									wire [12:0] b_imm = {instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
									// Trace: src/VX_decode.sv:34:5
									wire [20:0] jal_imm = {instr[31], instr[19:12], instr[20], instr[30:21], 1'b0};
									// Trace: src/VX_decode.sv:35:5
									reg [3:0] r_type;
									// Trace: src/VX_decode.sv:36:5
									always @(*)
										// Trace: src/VX_decode.sv:37:9
										case (func3)
											3'h0:
												// Trace: src/VX_decode.sv:38:19
												r_type = (opcode[5] && func7[5] ? 4'b0111 : 4'b0000);
											3'h1:
												// Trace: src/VX_decode.sv:39:19
												r_type = 4'b1111;
											3'h2:
												// Trace: src/VX_decode.sv:40:19
												r_type = 4'b0101;
											3'h3:
												// Trace: src/VX_decode.sv:41:19
												r_type = 4'b0100;
											3'h4:
												// Trace: src/VX_decode.sv:42:19
												r_type = 4'b1110;
											3'h5:
												// Trace: src/VX_decode.sv:43:19
												r_type = (func7[5] ? 4'b1001 : 4'b1000);
											3'h6:
												// Trace: src/VX_decode.sv:44:19
												r_type = 4'b1101;
											3'h7:
												// Trace: src/VX_decode.sv:45:19
												r_type = 4'b1100;
										endcase
									// Trace: src/VX_decode.sv:48:5
									reg [3:0] b_type;
									// Trace: src/VX_decode.sv:49:5
									always @(*)
										// Trace: src/VX_decode.sv:50:9
										case (func3)
											3'h0:
												// Trace: src/VX_decode.sv:51:19
												b_type = 4'b0000;
											3'h1:
												// Trace: src/VX_decode.sv:52:19
												b_type = 4'b0010;
											3'h4:
												// Trace: src/VX_decode.sv:53:19
												b_type = 4'b0101;
											3'h5:
												// Trace: src/VX_decode.sv:54:19
												b_type = 4'b0111;
											3'h6:
												// Trace: src/VX_decode.sv:55:19
												b_type = 4'b0100;
											3'h7:
												// Trace: src/VX_decode.sv:56:19
												b_type = 4'b0110;
											default:
												// Trace: src/VX_decode.sv:57:22
												b_type = 1'sbx;
										endcase
									// Trace: src/VX_decode.sv:60:5
									reg [3:0] s_type;
									// Trace: src/VX_decode.sv:61:5
									always @(*)
										// Trace: src/VX_decode.sv:62:9
										case (u_12)
											12'h000:
												// Trace: src/VX_decode.sv:63:22
												s_type = 4'b1010;
											12'h001:
												// Trace: src/VX_decode.sv:64:22
												s_type = 4'b1011;
											12'h002:
												// Trace: src/VX_decode.sv:65:22
												s_type = 4'b1100;
											12'h102:
												// Trace: src/VX_decode.sv:66:22
												s_type = 4'b1101;
											12'h302:
												// Trace: src/VX_decode.sv:67:22
												s_type = 4'b1110;
											default:
												// Trace: src/VX_decode.sv:68:22
												s_type = 1'sbx;
										endcase
									// Trace: src/VX_decode.sv:71:5
									reg [2:0] m_type;
									// Trace: src/VX_decode.sv:72:5
									always @(*)
										// Trace: src/VX_decode.sv:73:9
										case (func3)
											3'h0:
												// Trace: src/VX_decode.sv:74:19
												m_type = 3'b000;
											3'h1:
												// Trace: src/VX_decode.sv:75:19
												m_type = 3'b010;
											3'h2:
												// Trace: src/VX_decode.sv:76:19
												m_type = 3'b011;
											3'h3:
												// Trace: src/VX_decode.sv:77:19
												m_type = 3'b001;
											3'h4:
												// Trace: src/VX_decode.sv:78:19
												m_type = 3'b100;
											3'h5:
												// Trace: src/VX_decode.sv:79:19
												m_type = 3'b101;
											3'h6:
												// Trace: src/VX_decode.sv:80:19
												m_type = 3'b110;
											3'h7:
												// Trace: src/VX_decode.sv:81:19
												m_type = 3'b111;
										endcase
									// Trace: src/VX_decode.sv:89:5
									always @(*) begin
										// Trace: src/VX_decode.sv:90:9
										ex_type = 1'sbx;
										// Trace: src/VX_decode.sv:91:9
										op_type = 1'sbx;
										// Trace: src/VX_decode.sv:92:9
										op_args = 1'sbx;
										// Trace: src/VX_decode.sv:93:9
										rd_v = 1'sb0;
										// Trace: src/VX_decode.sv:94:9
										rs1_v = 1'sb0;
										// Trace: src/VX_decode.sv:95:9
										rs2_v = 1'sb0;
										// Trace: src/VX_decode.sv:96:9
										rs3_v = 1'sb0;
										// Trace: src/VX_decode.sv:97:9
										use_rd = 0;
										// Trace: src/VX_decode.sv:98:9
										use_rs1 = 0;
										// Trace: src/VX_decode.sv:99:9
										use_rs2 = 0;
										// Trace: src/VX_decode.sv:100:9
										use_rs3 = 0;
										// Trace: src/VX_decode.sv:101:9
										is_wstall = 0;
										// Trace: src/VX_decode.sv:102:9
										case (opcode)
											7'b0010011: begin
												// Trace: src/VX_decode.sv:104:17
												ex_type = 0;
												// Trace: src/VX_decode.sv:105:17
												op_type = r_type;
												// Trace: src/VX_decode.sv:106:17
												op_args[33-:2] = 0;
												// Trace: src/VX_decode.sv:107:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:108:17
												op_args[36] = 0;
												// Trace: src/VX_decode.sv:109:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:110:17
												op_args[31-:32] = {{21 {i_imm[11]}}, i_imm[10:0]};
												// Trace: src/VX_decode.sv:111:17
												use_rd = 1;
												// Trace: src/VX_decode.sv:112:9
												rd_v = {1'b0, rd};
												// Trace: src/VX_decode.sv:113:9
												use_rd = 1;
												// Trace: src/VX_decode.sv:114:9
												rs1_v = {1'b0, rs1};
												// Trace: src/VX_decode.sv:115:9
												use_rs1 = 1;
											end
											7'b0110011: begin
												// Trace: src/VX_decode.sv:118:17
												ex_type = 0;
												// Trace: src/VX_decode.sv:119:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:120:17
												op_args[36] = 0;
												// Trace: src/VX_decode.sv:121:17
												op_args[35] = 0;
												// Trace: src/VX_decode.sv:122:17
												use_rd = 1;
												// Trace: src/VX_decode.sv:123:9
												rd_v = {1'b0, rd};
												// Trace: src/VX_decode.sv:124:9
												use_rd = 1;
												// Trace: src/VX_decode.sv:125:9
												rs1_v = {1'b0, rs1};
												// Trace: src/VX_decode.sv:126:9
												use_rs1 = 1;
												// Trace: src/VX_decode.sv:127:9
												rs2_v = {1'b0, rs2};
												// Trace: src/VX_decode.sv:128:9
												use_rs2 = 1;
												// Trace: src/VX_decode.sv:129:17
												case (func7)
													7'b0000001: begin
														// Trace: src/VX_decode.sv:131:25
														op_type = sv2v_cast_4(m_type);
														// Trace: src/VX_decode.sv:132:25
														op_args[33-:2] = 2;
													end
													7'b0000111: begin
														// Trace: src/VX_decode.sv:135:25
														op_type = (func3[1] ? 4'b1011 : 4'b1010);
														// Trace: src/VX_decode.sv:136:25
														op_args[33-:2] = 0;
													end
													default: begin
														// Trace: src/VX_decode.sv:139:25
														op_type = r_type;
														// Trace: src/VX_decode.sv:140:25
														op_args[33-:2] = 0;
													end
												endcase
											end
											7'b0110111: begin
												// Trace: src/VX_decode.sv:145:17
												ex_type = 0;
												// Trace: src/VX_decode.sv:146:17
												op_type = 4'b0010;
												// Trace: src/VX_decode.sv:147:17
												op_args[33-:2] = 0;
												// Trace: src/VX_decode.sv:148:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:149:17
												op_args[36] = 0;
												// Trace: src/VX_decode.sv:150:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:151:17
												op_args[31-:32] = {ui_imm[19], ui_imm[18:0], 12'sd0};
												// Trace: src/VX_decode.sv:152:17
												use_rd = 1;
												// Trace: src/VX_decode.sv:153:9
												rd_v = {1'b0, rd};
												// Trace: src/VX_decode.sv:154:9
												use_rd = 1;
											end
											7'b0010111: begin
												// Trace: src/VX_decode.sv:157:17
												ex_type = 0;
												// Trace: src/VX_decode.sv:158:17
												op_type = 4'b0011;
												// Trace: src/VX_decode.sv:159:17
												op_args[33-:2] = 0;
												// Trace: src/VX_decode.sv:160:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:161:17
												op_args[36] = 1;
												// Trace: src/VX_decode.sv:162:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:163:17
												op_args[31-:32] = {ui_imm[19], ui_imm[18:0], 12'sd0};
												// Trace: src/VX_decode.sv:164:17
												use_rd = 1;
												// Trace: src/VX_decode.sv:165:9
												rd_v = {1'b0, rd};
												// Trace: src/VX_decode.sv:166:9
												use_rd = 1;
											end
											7'b1101111: begin
												// Trace: src/VX_decode.sv:169:17
												ex_type = 0;
												// Trace: src/VX_decode.sv:170:17
												op_type = 4'b1000;
												// Trace: src/VX_decode.sv:171:17
												op_args[33-:2] = 1;
												// Trace: src/VX_decode.sv:172:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:173:17
												op_args[36] = 1;
												// Trace: src/VX_decode.sv:174:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:175:17
												op_args[31-:32] = {{12 {jal_imm[20]}}, jal_imm[19:0]};
												// Trace: src/VX_decode.sv:176:17
												use_rd = 1;
												// Trace: src/VX_decode.sv:177:17
												is_wstall = 1;
												// Trace: src/VX_decode.sv:178:9
												rd_v = {1'b0, rd};
												// Trace: src/VX_decode.sv:179:9
												use_rd = 1;
											end
											7'b1100111: begin
												// Trace: src/VX_decode.sv:182:17
												ex_type = 0;
												// Trace: src/VX_decode.sv:183:17
												op_type = 4'b1001;
												// Trace: src/VX_decode.sv:184:17
												op_args[33-:2] = 1;
												// Trace: src/VX_decode.sv:185:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:186:17
												op_args[36] = 0;
												// Trace: src/VX_decode.sv:187:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:188:17
												op_args[31-:32] = {{21 {u_12[11]}}, u_12[10:0]};
												// Trace: src/VX_decode.sv:189:17
												use_rd = 1;
												// Trace: src/VX_decode.sv:190:17
												is_wstall = 1;
												// Trace: src/VX_decode.sv:191:9
												rd_v = {1'b0, rd};
												// Trace: src/VX_decode.sv:192:9
												use_rd = 1;
												// Trace: src/VX_decode.sv:193:9
												rs1_v = {1'b0, rs1};
												// Trace: src/VX_decode.sv:194:9
												use_rs1 = 1;
											end
											7'b1100011: begin
												// Trace: src/VX_decode.sv:197:17
												ex_type = 0;
												// Trace: src/VX_decode.sv:198:17
												op_type = b_type;
												// Trace: src/VX_decode.sv:199:17
												op_args[33-:2] = 1;
												// Trace: src/VX_decode.sv:200:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:201:17
												op_args[36] = 1;
												// Trace: src/VX_decode.sv:202:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:203:17
												op_args[31-:32] = {{20 {b_imm[12]}}, b_imm[11:0]};
												// Trace: src/VX_decode.sv:204:17
												is_wstall = 1;
												// Trace: src/VX_decode.sv:205:9
												rs1_v = {1'b0, rs1};
												// Trace: src/VX_decode.sv:206:9
												use_rs1 = 1;
												// Trace: src/VX_decode.sv:207:9
												rs2_v = {1'b0, rs2};
												// Trace: src/VX_decode.sv:208:9
												use_rs2 = 1;
											end
											7'b0001111: begin
												// Trace: src/VX_decode.sv:211:17
												ex_type = 1;
												// Trace: src/VX_decode.sv:212:17
												op_type = 4'b1111;
												// Trace: src/VX_decode.sv:213:17
												op_args[13] = 0;
												// Trace: src/VX_decode.sv:214:17
												op_args[12] = 0;
												// Trace: src/VX_decode.sv:215:17
												op_args[11-:12] = 0;
											end
											7'b1110011:
												// Trace: src/VX_decode.sv:218:17
												if (func3[1:0] != 0) begin
													// Trace: src/VX_decode.sv:219:21
													ex_type = 2;
													// Trace: src/VX_decode.sv:220:21
													op_type = sv2v_cast_4((4'h6 + sv2v_cast_4(func3[1:0])) - 4'h1);
													// Trace: src/VX_decode.sv:221:21
													op_args[16-:12] = u_12;
													// Trace: src/VX_decode.sv:222:21
													op_args[17] = func3[2];
													// Trace: src/VX_decode.sv:223:21
													use_rd = 1;
													// Trace: src/VX_decode.sv:224:21
													is_wstall = is_fpu_csr;
													// Trace: src/VX_decode.sv:225:9
													rd_v = {1'b0, rd};
													// Trace: src/VX_decode.sv:226:9
													use_rd = 1;
													// Trace: src/VX_decode.sv:227:21
													if (func3[2])
														// Trace: src/VX_decode.sv:228:25
														op_args[4-:5] = rs1;
													else begin
														// Trace: src/VX_decode.sv:230:9
														rs1_v = {1'b0, rs1};
														// Trace: src/VX_decode.sv:231:9
														use_rs1 = 1;
													end
												end
												else begin
													// Trace: src/VX_decode.sv:234:21
													ex_type = 0;
													// Trace: src/VX_decode.sv:235:21
													op_type = s_type;
													// Trace: src/VX_decode.sv:236:21
													op_args[33-:2] = 1;
													// Trace: src/VX_decode.sv:237:21
													op_args[34] = 0;
													// Trace: src/VX_decode.sv:238:21
													op_args[35] = 1;
													// Trace: src/VX_decode.sv:239:21
													op_args[36] = 1;
													// Trace: src/VX_decode.sv:240:21
													op_args[31-:32] = 32'd4;
													// Trace: src/VX_decode.sv:241:21
													use_rd = 1;
													// Trace: src/VX_decode.sv:242:21
													is_wstall = 1;
													// Trace: src/VX_decode.sv:243:9
													rd_v = {1'b0, rd};
													// Trace: src/VX_decode.sv:244:9
													use_rd = 1;
												end
											7'b0000111, 7'b0000011: begin
												// Trace: src/VX_decode.sv:249:17
												ex_type = 1;
												// Trace: src/VX_decode.sv:250:17
												op_type = sv2v_cast_4({1'b0, func3});
												// Trace: src/VX_decode.sv:251:17
												op_args[13] = 0;
												// Trace: src/VX_decode.sv:252:17
												op_args[12] = opcode[2];
												// Trace: src/VX_decode.sv:253:17
												op_args[11-:12] = u_12;
												// Trace: src/VX_decode.sv:254:17
												use_rd = 1;
												// Trace: src/VX_decode.sv:255:17
												if (opcode[2]) begin
													// Trace: src/VX_decode.sv:256:9
													rd_v = {1'b1, rd};
													// Trace: src/VX_decode.sv:257:9
													use_rd = 1;
												end
												else
													// Trace: src/VX_decode.sv:259:9
													rd_v = {1'b0, rd};
												// Trace: src/VX_decode.sv:260:9
												use_rd = 1;
												// Trace: src/VX_decode.sv:261:9
												rs1_v = {1'b0, rs1};
												// Trace: src/VX_decode.sv:262:9
												use_rs1 = 1;
											end
											7'b0100111, 7'b0100011: begin
												// Trace: src/VX_decode.sv:266:17
												ex_type = 1;
												// Trace: src/VX_decode.sv:267:17
												op_type = sv2v_cast_4({1'b1, func3});
												// Trace: src/VX_decode.sv:268:17
												op_args[13] = 1;
												// Trace: src/VX_decode.sv:269:17
												op_args[12] = opcode[2];
												// Trace: src/VX_decode.sv:270:17
												op_args[11-:12] = s_imm;
												// Trace: src/VX_decode.sv:271:9
												rs1_v = {1'b0, rs1};
												// Trace: src/VX_decode.sv:272:9
												use_rs1 = 1;
												// Trace: src/VX_decode.sv:273:17
												if (opcode[2]) begin
													// Trace: src/VX_decode.sv:274:9
													rs2_v = {1'b1, rs2};
													// Trace: src/VX_decode.sv:275:9
													use_rs2 = 1;
												end
												else
													// Trace: src/VX_decode.sv:277:9
													rs2_v = {1'b0, rs2};
												// Trace: src/VX_decode.sv:278:9
												use_rs2 = 1;
											end
											7'b1000011, 7'b1000111, 7'b1001011, 7'b1001111: begin
												// Trace: src/VX_decode.sv:285:17
												ex_type = 3;
												// Trace: src/VX_decode.sv:286:17
												op_type = sv2v_cast_4({3'b001, opcode[3]});
												// Trace: src/VX_decode.sv:287:17
												op_args[4-:3] = func3;
												// Trace: src/VX_decode.sv:288:17
												op_args[0] = func2[0];
												// Trace: src/VX_decode.sv:289:17
												op_args[1] = opcode[3] ^ opcode[2];
												// Trace: src/VX_decode.sv:290:17
												use_rd = 1;
												// Trace: src/VX_decode.sv:291:9
												rd_v = {1'b1, rd};
												// Trace: src/VX_decode.sv:292:9
												use_rd = 1;
												// Trace: src/VX_decode.sv:293:9
												rs1_v = {1'b1, rs1};
												// Trace: src/VX_decode.sv:294:9
												use_rs1 = 1;
												// Trace: src/VX_decode.sv:295:9
												rs2_v = {1'b1, rs2};
												// Trace: src/VX_decode.sv:296:9
												use_rs2 = 1;
												// Trace: src/VX_decode.sv:297:9
												rs3_v = {1'b1, rs3};
												// Trace: src/VX_decode.sv:298:9
												use_rs3 = 1;
											end
											7'b1010011: begin
												// Trace: src/VX_decode.sv:301:17
												ex_type = 3;
												// Trace: src/VX_decode.sv:302:17
												op_args[4-:3] = func3;
												// Trace: src/VX_decode.sv:303:17
												op_args[0] = func2[0];
												// Trace: src/VX_decode.sv:304:17
												op_args[1] = rs2[1];
												// Trace: src/VX_decode.sv:305:17
												use_rd = 1;
												// Trace: src/VX_decode.sv:306:17
												case (func5)
													5'b00000, 5'b00001, 5'b00010: begin
														// Trace: src/VX_decode.sv:311:25
														op_type = sv2v_cast_4({3'b000, func5[1]});
														// Trace: src/VX_decode.sv:312:25
														op_args[1] = func5[0];
														// Trace: src/VX_decode.sv:313:9
														rd_v = {1'b1, rd};
														// Trace: src/VX_decode.sv:314:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:315:9
														rs1_v = {1'b1, rs1};
														// Trace: src/VX_decode.sv:316:9
														use_rs1 = 1;
														// Trace: src/VX_decode.sv:317:9
														rs2_v = {1'b1, rs2};
														// Trace: src/VX_decode.sv:318:9
														use_rs2 = 1;
													end
													5'b00100: begin
														// Trace: src/VX_decode.sv:321:25
														op_type = 4'b1110;
														// Trace: src/VX_decode.sv:322:25
														op_args[4-:3] = sv2v_cast_3(func3[1:0]);
														// Trace: src/VX_decode.sv:323:9
														rd_v = {1'b1, rd};
														// Trace: src/VX_decode.sv:324:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:325:9
														rs1_v = {1'b1, rs1};
														// Trace: src/VX_decode.sv:326:9
														use_rs1 = 1;
														// Trace: src/VX_decode.sv:327:9
														rs2_v = {1'b1, rs2};
														// Trace: src/VX_decode.sv:328:9
														use_rs2 = 1;
													end
													5'b00101: begin
														// Trace: src/VX_decode.sv:331:25
														op_type = 4'b1110;
														// Trace: src/VX_decode.sv:332:25
														op_args[4-:3] = sv2v_cast_3_signed((func3[0] ? 7 : 6));
														// Trace: src/VX_decode.sv:333:9
														rd_v = {1'b1, rd};
														// Trace: src/VX_decode.sv:334:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:335:9
														rs1_v = {1'b1, rs1};
														// Trace: src/VX_decode.sv:336:9
														use_rs1 = 1;
														// Trace: src/VX_decode.sv:337:9
														rs2_v = {1'b1, rs2};
														// Trace: src/VX_decode.sv:338:9
														use_rs2 = 1;
													end
													5'b00011: begin
														// Trace: src/VX_decode.sv:341:25
														op_type = 4'b0100;
														// Trace: src/VX_decode.sv:342:9
														rd_v = {1'b1, rd};
														// Trace: src/VX_decode.sv:343:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:344:9
														rs1_v = {1'b1, rs1};
														// Trace: src/VX_decode.sv:345:9
														use_rs1 = 1;
														// Trace: src/VX_decode.sv:346:9
														rs2_v = {1'b1, rs2};
														// Trace: src/VX_decode.sv:347:9
														use_rs2 = 1;
													end
													5'b01011: begin
														// Trace: src/VX_decode.sv:350:25
														op_type = 4'b0101;
														// Trace: src/VX_decode.sv:351:9
														rd_v = {1'b1, rd};
														// Trace: src/VX_decode.sv:352:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:353:9
														rs1_v = {1'b1, rs1};
														// Trace: src/VX_decode.sv:354:9
														use_rs1 = 1;
													end
													5'b10100: begin
														// Trace: src/VX_decode.sv:357:25
														op_type = 4'b1100;
														// Trace: src/VX_decode.sv:358:9
														rd_v = {1'b0, rd};
														// Trace: src/VX_decode.sv:359:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:360:9
														rs1_v = {1'b1, rs1};
														// Trace: src/VX_decode.sv:361:9
														use_rs1 = 1;
														// Trace: src/VX_decode.sv:362:9
														rs2_v = {1'b1, rs2};
														// Trace: src/VX_decode.sv:363:9
														use_rs2 = 1;
													end
													5'b11000: begin
														// Trace: src/VX_decode.sv:366:25
														op_type = (rs2[0] ? 4'b1001 : 4'b1000);
														// Trace: src/VX_decode.sv:367:9
														rd_v = {1'b0, rd};
														// Trace: src/VX_decode.sv:368:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:369:9
														rs1_v = {1'b1, rs1};
														// Trace: src/VX_decode.sv:370:9
														use_rs1 = 1;
													end
													5'b11010: begin
														// Trace: src/VX_decode.sv:373:25
														op_type = (rs2[0] ? 4'b1011 : 4'b1010);
														// Trace: src/VX_decode.sv:374:9
														rd_v = {1'b1, rd};
														// Trace: src/VX_decode.sv:375:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:376:9
														rs1_v = {1'b0, rs1};
														// Trace: src/VX_decode.sv:377:9
														use_rs1 = 1;
													end
													5'b11100: begin
														// Trace: src/VX_decode.sv:380:25
														if (func3[0]) begin
															// Trace: src/VX_decode.sv:381:29
															op_type = 4'b1110;
															// Trace: src/VX_decode.sv:382:29
															op_args[4-:3] = 3'sd3;
														end
														else begin
															// Trace: src/VX_decode.sv:384:29
															op_type = 4'b1110;
															// Trace: src/VX_decode.sv:385:29
															op_args[4-:3] = 3'sd4;
														end
														// Trace: src/VX_decode.sv:387:9
														rd_v = {1'b0, rd};
														// Trace: src/VX_decode.sv:388:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:389:9
														rs1_v = {1'b1, rs1};
														// Trace: src/VX_decode.sv:390:9
														use_rs1 = 1;
													end
													5'b11110: begin
														// Trace: src/VX_decode.sv:393:25
														op_type = 4'b1110;
														// Trace: src/VX_decode.sv:394:25
														op_args[4-:3] = 3'sd5;
														// Trace: src/VX_decode.sv:395:9
														rd_v = {1'b1, rd};
														// Trace: src/VX_decode.sv:396:9
														use_rd = 1;
														// Trace: src/VX_decode.sv:397:9
														rs1_v = {1'b0, rs1};
														// Trace: src/VX_decode.sv:398:9
														use_rs1 = 1;
													end
													default:
														;
												endcase
											end
											7'b0001011:
												// Trace: src/VX_decode.sv:404:17
												case (func7)
													7'h00: begin
														// Trace: src/VX_decode.sv:406:25
														ex_type = 2;
														// Trace: src/VX_decode.sv:407:25
														is_wstall = 1;
														// Trace: src/VX_decode.sv:408:25
														case (func3)
															3'h0: begin
																// Trace: src/VX_decode.sv:410:33
																op_type = 4'h0;
																// Trace: src/VX_decode.sv:411:9
																rs1_v = {1'b0, rs1};
																// Trace: src/VX_decode.sv:412:9
																use_rs1 = 1;
															end
															3'h1: begin
																// Trace: src/VX_decode.sv:415:33
																op_type = 4'h1;
																// Trace: src/VX_decode.sv:416:9
																rs1_v = {1'b0, rs1};
																// Trace: src/VX_decode.sv:417:9
																use_rs1 = 1;
																// Trace: src/VX_decode.sv:418:9
																rs2_v = {1'b0, rs2};
																// Trace: src/VX_decode.sv:419:9
																use_rs2 = 1;
															end
															3'h2: begin
																// Trace: src/VX_decode.sv:422:33
																op_type = 4'h2;
																// Trace: src/VX_decode.sv:423:33
																use_rd = 1;
																// Trace: src/VX_decode.sv:424:33
																op_args[0] = rs2[0];
																// Trace: src/VX_decode.sv:425:9
																rs1_v = {1'b0, rs1};
																// Trace: src/VX_decode.sv:426:9
																use_rs1 = 1;
																// Trace: src/VX_decode.sv:427:9
																rd_v = {1'b0, rd};
																// Trace: src/VX_decode.sv:428:9
																use_rd = 1;
															end
															3'h3: begin
																// Trace: src/VX_decode.sv:431:33
																op_type = 4'h3;
																// Trace: src/VX_decode.sv:432:9
																rs1_v = {1'b0, rs1};
																// Trace: src/VX_decode.sv:433:9
																use_rs1 = 1;
															end
															3'h4: begin
																// Trace: src/VX_decode.sv:436:33
																op_type = 4'h4;
																// Trace: src/VX_decode.sv:437:9
																rs1_v = {1'b0, rs1};
																// Trace: src/VX_decode.sv:438:9
																use_rs1 = 1;
																// Trace: src/VX_decode.sv:439:9
																rs2_v = {1'b0, rs2};
																// Trace: src/VX_decode.sv:440:9
																use_rs2 = 1;
															end
															3'h5: begin
																// Trace: src/VX_decode.sv:443:33
																op_type = 4'h5;
																// Trace: src/VX_decode.sv:444:33
																op_args[0] = rd[0];
																// Trace: src/VX_decode.sv:445:9
																rs1_v = {1'b0, rs1};
																// Trace: src/VX_decode.sv:446:9
																use_rs1 = 1;
																// Trace: src/VX_decode.sv:447:9
																rs2_v = {1'b0, rs2};
																// Trace: src/VX_decode.sv:448:9
																use_rs2 = 1;
															end
															default:
																;
														endcase
													end
													default:
														;
												endcase
											default:
												;
										endcase
									end
									// Trace: src/VX_decode.sv:459:5
									wire wb = use_rd && (rd_v != 0);
									// Trace: src/VX_decode.sv:460:5
									VX_elastic_buffer #(
										.DATAW(DATAW),
										.SIZE(0)
									) req_buf(
										.clk(clk),
										.reset(reset),
										.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.valid),
										.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.ready),
										.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[69], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[68-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[66-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[62-:31], ex_type, op_type, op_args, wb, rd_v, rs1_v, rs2_v, rs3_v}),
										.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[105], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[104-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[102-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[98-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[67-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[65-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[61-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[24], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[23-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[17-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[11-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[5-:6]}),
										.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.valid),
										.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.ready)
									);
									// Trace: src/VX_decode.sv:473:5
									wire fetch_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.ready;
									// Trace: src/VX_decode.sv:474:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.valid = fetch_fire;
									// Trace: src/VX_decode.sv:475:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[68-:2];
									// Trace: src/VX_decode.sv:476:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.unlock = ~is_wstall;
								end
								assign decode.clk = clk;
								assign decode.reset = reset;
								// Trace: src/VX_core.sv:70:5
								// expanded module instance: issue
								localparam _bbase_CF65A_writeback_if = 0;
								localparam _bbase_CF65A_dispatch_if = 0;
								localparam _param_CF65A_INSTANCE_ID = "";
								if (1) begin : issue
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_issue.sv:2:16
									localparam INSTANCE_ID = _param_CF65A_INSTANCE_ID;
									// Trace: src/VX_issue.sv:4:5
									wire clk;
									// Trace: src/VX_issue.sv:5:5
									wire reset;
									// Trace: src/VX_issue.sv:6:5
									// removed modport instance decode_if
									// Trace: src/VX_issue.sv:7:5
									localparam _mbase_writeback_if = 0;
									// Trace: src/VX_issue.sv:8:5
									localparam _mbase_dispatch_if = 0;
									// Trace: src/VX_issue.sv:10:5
									localparam VX_gpu_pkg_ISSUE_ISW = 0;
									localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
									function [0:0] VX_gpu_pkg_wid_to_isw;
										// Trace: src/VX_gpu_pkg.sv:163:9
										input reg [1:0] wid;
										// Trace: src/VX_gpu_pkg.sv:165:9
										begin
											// Trace: src/VX_gpu_pkg.sv:168:13
											VX_gpu_pkg_wid_to_isw = 0;
										end
									endfunction
									wire [0:0] decode_isw = VX_gpu_pkg_wid_to_isw(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[104-:2]);
									// Trace: src/VX_issue.sv:11:5
									localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
									localparam VX_gpu_pkg_ISSUE_WIS = 2;
									localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
									function [1:0] VX_gpu_pkg_wid_to_wis;
										// Trace: src/VX_gpu_pkg.sv:172:9
										input reg [1:0] wid;
										// Trace: src/VX_gpu_pkg.sv:174:9
										begin
											// Trace: src/VX_gpu_pkg.sv:175:13
											VX_gpu_pkg_wid_to_wis = wid >> VX_gpu_pkg_ISSUE_ISW;
										end
									endfunction
									wire [1:0] decode_wis = VX_gpu_pkg_wid_to_wis(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[104-:2]);
									// Trace: src/VX_issue.sv:12:5
									wire [0:0] decode_ready_in;
									// Trace: src/VX_issue.sv:13:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.ready = decode_ready_in[decode_isw];
									// Trace: src/VX_issue.sv:15:5
									genvar _gv_issue_id_1;
									for (_gv_issue_id_1 = 0; _gv_issue_id_1 < 1; _gv_issue_id_1 = _gv_issue_id_1 + 1) begin : g_slices
										localparam issue_id = _gv_issue_id_1;
										// Trace: src/VX_issue.sv:16:9
										// expanded interface instance: per_issue_decode_if
										localparam _param_5C540_NUM_WARPS = VX_gpu_pkg_PER_ISSUE_WARPS;
										if (1) begin : per_issue_decode_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_decode_if.sv:2:15
											localparam NUM_WARPS = _param_5C540_NUM_WARPS;
											// Trace: src/VX_decode_if.sv:3:15
											localparam NW_WIDTH = 2;
											// Trace: src/VX_decode_if.sv:5:5
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_decode_if.sv:19:5
											wire valid;
											// Trace: src/VX_decode_if.sv:20:5
											wire [105:0] data;
											// Trace: src/VX_decode_if.sv:21:5
											wire ready;
											// Trace: src/VX_decode_if.sv:22:5
											// Trace: src/VX_decode_if.sv:27:5
										end
										// Trace: src/VX_issue.sv:19:9
										// expanded interface instance: per_issue_dispatch_if
										genvar _arr_18544;
										for (_arr_18544 = 0; _arr_18544 <= 3; _arr_18544 = _arr_18544 + 1) begin : per_issue_dispatch_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_dispatch_if.sv:2:5
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											localparam VX_gpu_pkg_ISSUE_WIS = 2;
											localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_dispatch_if.sv:16:5
											wire valid;
											// Trace: src/VX_dispatch_if.sv:17:5
											wire [471:0] data;
											// Trace: src/VX_dispatch_if.sv:18:5
											wire ready;
											// Trace: src/VX_dispatch_if.sv:19:5
											// Trace: src/VX_dispatch_if.sv:24:5
										end
										// Trace: src/VX_issue.sv:20:9
										assign per_issue_decode_if.valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.valid && (decode_isw == sv2v_cast_1_signed(issue_id));
										// Trace: src/VX_issue.sv:21:9
										assign per_issue_decode_if.data[105] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[105];
										// Trace: src/VX_issue.sv:22:9
										assign per_issue_decode_if.data[104-:2] = decode_wis;
										// Trace: src/VX_issue.sv:23:9
										assign per_issue_decode_if.data[102-:4] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[102-:4];
										// Trace: src/VX_issue.sv:24:9
										assign per_issue_decode_if.data[98-:31] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[98-:31];
										// Trace: src/VX_issue.sv:25:9
										assign per_issue_decode_if.data[67-:2] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[67-:2];
										// Trace: src/VX_issue.sv:26:9
										assign per_issue_decode_if.data[65-:4] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[65-:4];
										// Trace: src/VX_issue.sv:27:9
										assign per_issue_decode_if.data[61-:37] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[61-:37];
										// Trace: src/VX_issue.sv:28:9
										assign per_issue_decode_if.data[24] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[24];
										// Trace: src/VX_issue.sv:29:9
										assign per_issue_decode_if.data[23-:6] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[23-:6];
										// Trace: src/VX_issue.sv:30:9
										assign per_issue_decode_if.data[17-:6] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[17-:6];
										// Trace: src/VX_issue.sv:31:9
										assign per_issue_decode_if.data[11-:6] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[11-:6];
										// Trace: src/VX_issue.sv:32:9
										assign per_issue_decode_if.data[5-:6] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[5-:6];
										// Trace: src/VX_issue.sv:33:9
										assign decode_ready_in[issue_id] = per_issue_decode_if.ready;
										// Trace: src/VX_issue.sv:34:9
										// expanded module instance: issue_slice
										localparam _bbase_A8822_writeback_if = issue_id + _mbase_writeback_if;
										localparam _bbase_A8822_dispatch_if = 0;
										localparam _param_A8822_INSTANCE_ID = "";
										localparam _param_A8822_ISSUE_ID = issue_id;
										if (1) begin : issue_slice
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_issue_slice.sv:2:16
											localparam INSTANCE_ID = _param_A8822_INSTANCE_ID;
											// Trace: src/VX_issue_slice.sv:3:15
											localparam ISSUE_ID = _param_A8822_ISSUE_ID;
											// Trace: src/VX_issue_slice.sv:5:5
											wire clk;
											// Trace: src/VX_issue_slice.sv:6:5
											wire reset;
											// Trace: src/VX_issue_slice.sv:7:5
											// removed modport instance decode_if
											// Trace: src/VX_issue_slice.sv:8:5
											localparam _mbase_writeback_if = _bbase_A8822_writeback_if;
											// Trace: src/VX_issue_slice.sv:9:5
											localparam _mbase_dispatch_if = 0;
											// Trace: src/VX_issue_slice.sv:11:5
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											// expanded interface instance: ibuffer_if
											genvar _arr_F0EBA;
											for (_arr_F0EBA = 0; _arr_F0EBA <= 3; _arr_F0EBA = _arr_F0EBA + 1) begin : ibuffer_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_ibuffer_if.sv:2:5
												// removed localparam type VX_gpu_pkg_alu_args_t
												// removed localparam type VX_gpu_pkg_csr_args_t
												// removed localparam type VX_gpu_pkg_fpu_args_t
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												// removed localparam type data_t
												// Trace: src/VX_ibuffer_if.sv:15:5
												wire valid;
												// Trace: src/VX_ibuffer_if.sv:16:5
												wire [103:0] data;
												// Trace: src/VX_ibuffer_if.sv:17:5
												wire ready;
												// Trace: src/VX_ibuffer_if.sv:18:5
												// Trace: src/VX_ibuffer_if.sv:23:5
											end
											// Trace: src/VX_issue_slice.sv:12:5
											// expanded interface instance: scoreboard_if
											if (1) begin : scoreboard_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_scoreboard_if.sv:2:5
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam VX_gpu_pkg_ISSUE_WIS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
												// removed localparam type VX_gpu_pkg_alu_args_t
												// removed localparam type VX_gpu_pkg_csr_args_t
												// removed localparam type VX_gpu_pkg_fpu_args_t
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												// removed localparam type data_t
												// Trace: src/VX_scoreboard_if.sv:16:5
												wire valid;
												// Trace: src/VX_scoreboard_if.sv:17:5
												wire [105:0] data;
												// Trace: src/VX_scoreboard_if.sv:18:5
												wire ready;
												// Trace: src/VX_scoreboard_if.sv:19:5
												// Trace: src/VX_scoreboard_if.sv:24:5
											end
											// Trace: src/VX_issue_slice.sv:13:5
											// expanded interface instance: operands_if
											if (1) begin : operands_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_operands_if.sv:2:5
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam VX_gpu_pkg_ISSUE_WIS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
												// removed localparam type VX_gpu_pkg_alu_args_t
												// removed localparam type VX_gpu_pkg_csr_args_t
												// removed localparam type VX_gpu_pkg_fpu_args_t
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												// removed localparam type data_t
												// Trace: src/VX_operands_if.sv:16:5
												wire valid;
												// Trace: src/VX_operands_if.sv:17:5
												wire [471:0] data;
												// Trace: src/VX_operands_if.sv:18:5
												wire ready;
												// Trace: src/VX_operands_if.sv:19:5
												// Trace: src/VX_operands_if.sv:24:5
											end
											// Trace: src/VX_issue_slice.sv:14:5
											// expanded module instance: ibuffer
											localparam _bbase_D579A_ibuffer_if = 0;
											localparam _param_D579A_INSTANCE_ID = "";
											if (1) begin : ibuffer
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_ibuffer.sv:2:16
												localparam INSTANCE_ID = _param_D579A_INSTANCE_ID;
												// Trace: src/VX_ibuffer.sv:4:5
												wire clk;
												// Trace: src/VX_ibuffer.sv:5:5
												wire reset;
												// Trace: src/VX_ibuffer.sv:6:5
												// removed modport instance decode_if
												// Trace: src/VX_ibuffer.sv:7:5
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam _mbase_ibuffer_if = 0;
												// Trace: src/VX_ibuffer.sv:9:5
												// removed localparam type VX_gpu_pkg_alu_args_t
												// removed localparam type VX_gpu_pkg_csr_args_t
												// removed localparam type VX_gpu_pkg_fpu_args_t
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam DATAW = 104;
												// Trace: src/VX_ibuffer.sv:10:5
												wire [3:0] ibuf_ready_in;
												// Trace: src/VX_ibuffer.sv:11:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.ready = ibuf_ready_in[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[104-:2]];
												// Trace: src/VX_ibuffer.sv:12:5
												genvar _gv_w_1;
												localparam VX_gpu_pkg_ISSUE_WIS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
												for (_gv_w_1 = 0; _gv_w_1 < VX_gpu_pkg_PER_ISSUE_WARPS; _gv_w_1 = _gv_w_1 + 1) begin : g_instr_bufs
													localparam w = _gv_w_1;
													// Trace: src/VX_ibuffer.sv:13:9
													VX_elastic_buffer #(
														.DATAW(DATAW),
														.SIZE(4),
														.OUT_REG(1)
													) instr_buf(
														.clk(clk),
														.reset(reset),
														.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.valid && (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[104-:2] == sv2v_cast_2_signed(w))),
														.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[105], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[102-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[98-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[67-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[65-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[61-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[24], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[23-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[17-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[11-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_decode_if.data[5-:6]}),
														.ready_in(ibuf_ready_in[w]),
														.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].valid),
														.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data),
														.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].ready)
													);
												end
											end
											assign ibuffer.clk = clk;
											assign ibuffer.reset = reset;
											// Trace: src/VX_issue_slice.sv:22:5
											// expanded module instance: scoreboard
											localparam _bbase_85D2C_writeback_if = issue_id + _mbase_writeback_if;
											localparam _bbase_85D2C_ibuffer_if = 0;
											localparam _param_85D2C_INSTANCE_ID = "";
											if (1) begin : scoreboard
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_scoreboard.sv:2:16
												localparam INSTANCE_ID = _param_85D2C_INSTANCE_ID;
												// Trace: src/VX_scoreboard.sv:4:5
												wire clk;
												// Trace: src/VX_scoreboard.sv:5:5
												wire reset;
												// Trace: src/VX_scoreboard.sv:6:5
												localparam _mbase_writeback_if = _bbase_85D2C_writeback_if;
												// Trace: src/VX_scoreboard.sv:7:5
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam _mbase_ibuffer_if = 0;
												// Trace: src/VX_scoreboard.sv:8:5
												// removed modport instance scoreboard_if
												// Trace: src/VX_scoreboard.sv:10:5
												localparam NUM_SRC_OPDS = 3;
												// Trace: src/VX_scoreboard.sv:11:5
												localparam NUM_OPDS = 4;
												// Trace: src/VX_scoreboard.sv:12:5
												// removed localparam type VX_gpu_pkg_alu_args_t
												// removed localparam type VX_gpu_pkg_csr_args_t
												// removed localparam type VX_gpu_pkg_fpu_args_t
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam DATAW = 104;
												// Trace: src/VX_scoreboard.sv:13:5
												// expanded interface instance: staging_if
												genvar _arr_8EA22;
												for (_arr_8EA22 = 0; _arr_8EA22 <= 3; _arr_8EA22 = _arr_8EA22 + 1) begin : staging_if
													// removed import VX_gpu_pkg::*;
													// Trace: src/VX_ibuffer_if.sv:2:5
													// removed localparam type VX_gpu_pkg_alu_args_t
													// removed localparam type VX_gpu_pkg_csr_args_t
													// removed localparam type VX_gpu_pkg_fpu_args_t
													// removed localparam type VX_gpu_pkg_lsu_args_t
													// removed localparam type VX_gpu_pkg_wctl_args_t
													// removed localparam type VX_gpu_pkg_op_args_t
													// removed localparam type data_t
													// Trace: src/VX_ibuffer_if.sv:15:5
													wire valid;
													// Trace: src/VX_ibuffer_if.sv:16:5
													wire [103:0] data;
													// Trace: src/VX_ibuffer_if.sv:17:5
													wire ready;
													// Trace: src/VX_ibuffer_if.sv:18:5
													// Trace: src/VX_ibuffer_if.sv:23:5
												end
												// Trace: src/VX_scoreboard.sv:14:5
												reg [3:0] operands_ready;
												// Trace: src/VX_scoreboard.sv:15:5
												genvar _gv_w_2;
												for (_gv_w_2 = 0; _gv_w_2 < VX_gpu_pkg_PER_ISSUE_WARPS; _gv_w_2 = _gv_w_2 + 1) begin : g_stanging_bufs
													localparam w = _gv_w_2;
													// Trace: src/VX_scoreboard.sv:16:9
													VX_pipe_buffer #(.DATAW(DATAW)) stanging_buf(
														.clk(clk),
														.reset(reset),
														.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].valid),
														.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data),
														.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].ready),
														.valid_out(staging_if[w].valid),
														.data_out(staging_if[w].data),
														.ready_out(staging_if[w].ready)
													);
												end
												// Trace: src/VX_scoreboard.sv:29:5
												genvar _gv_w_3;
												localparam VX_gpu_pkg_ISSUE_WIS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
												for (_gv_w_3 = 0; _gv_w_3 < VX_gpu_pkg_PER_ISSUE_WARPS; _gv_w_3 = _gv_w_3 + 1) begin : g_scoreboard
													localparam w = _gv_w_3;
													// Trace: src/VX_scoreboard.sv:30:9
													reg [63:0] inuse_regs;
													// Trace: src/VX_scoreboard.sv:31:9
													reg [3:0] operands_busy;
													reg [3:0] operands_busy_n;
													// Trace: src/VX_scoreboard.sv:32:9
													wire ibuffer_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].ready;
													// Trace: src/VX_scoreboard.sv:33:9
													wire staging_fire = staging_if[w].valid && staging_if[w].ready;
													// Trace: src/VX_scoreboard.sv:34:9
													wire writeback_fire = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].valid && (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[172-:2] == sv2v_cast_2_signed(w))) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[0];
													// Trace: src/VX_scoreboard.sv:37:9
													wire [23:0] ibuf_opds;
													wire [23:0] stg_opds;
													// Trace: src/VX_scoreboard.sv:38:9
													assign ibuf_opds = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[5-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[11-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[17-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[23-:6]};
													// Trace: src/VX_scoreboard.sv:39:9
													assign stg_opds = {staging_if[w].data[5-:6], staging_if[w].data[11-:6], staging_if[w].data[17-:6], staging_if[w].data[23-:6]};
													// Trace: src/VX_scoreboard.sv:40:9
													always @(*)
														// Trace: src/VX_scoreboard.sv:41:13
														begin : sv2v_autoblock_5
															// Trace: src/VX_scoreboard.sv:41:18
															integer i;
															// Trace: src/VX_scoreboard.sv:41:18
															for (i = 0; i < NUM_OPDS; i = i + 1)
																begin
																	// Trace: src/VX_scoreboard.sv:42:17
																	operands_busy_n[i] = operands_busy[i];
																	// Trace: src/VX_scoreboard.sv:43:17
																	if (ibuffer_fire)
																		// Trace: src/VX_scoreboard.sv:44:21
																		operands_busy_n[i] = inuse_regs[ibuf_opds[i * 6+:6]];
																	if (writeback_fire) begin
																		begin
																			// Trace: src/VX_scoreboard.sv:47:21
																			if (ibuffer_fire) begin
																				begin
																					// Trace: src/VX_scoreboard.sv:48:25
																					if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[135-:6] == ibuf_opds[i * 6+:6])
																						// Trace: src/VX_scoreboard.sv:49:29
																						operands_busy_n[i] = 0;
																				end
																			end
																			else
																				// Trace: src/VX_scoreboard.sv:52:25
																				if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[135-:6] == stg_opds[i * 6+:6])
																					// Trace: src/VX_scoreboard.sv:53:29
																					operands_busy_n[i] = 0;
																		end
																	end
																	if ((staging_fire && staging_if[w].data[24]) && (staging_if[w].data[23-:6] == ibuf_opds[i * 6+:6]))
																		// Trace: src/VX_scoreboard.sv:58:21
																		operands_busy_n[i] = 1;
																end
														end
													// Trace: src/VX_scoreboard.sv:62:9
													always @(posedge clk) begin
														// Trace: src/VX_scoreboard.sv:63:13
														if (reset)
															// Trace: src/VX_scoreboard.sv:64:17
															inuse_regs <= 1'sb0;
														else begin
															// Trace: src/VX_scoreboard.sv:66:17
															if (writeback_fire)
																// Trace: src/VX_scoreboard.sv:67:21
																inuse_regs[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[135-:6]] <= 0;
															if (staging_fire && staging_if[w].data[24])
																// Trace: src/VX_scoreboard.sv:70:21
																inuse_regs[staging_if[w].data[23-:6]] <= 1;
														end
														// Trace: src/VX_scoreboard.sv:73:13
														operands_busy <= operands_busy_n;
														// Trace: src/VX_scoreboard.sv:74:13
														operands_ready[w] <= ~(|operands_busy_n);
													end
												end
												// Trace: src/VX_scoreboard.sv:77:5
												wire [3:0] arb_valid_in;
												// Trace: src/VX_scoreboard.sv:78:5
												wire [415:0] arb_data_in;
												// Trace: src/VX_scoreboard.sv:79:5
												wire [3:0] arb_ready_in;
												// Trace: src/VX_scoreboard.sv:80:5
												genvar _gv_w_4;
												for (_gv_w_4 = 0; _gv_w_4 < VX_gpu_pkg_PER_ISSUE_WARPS; _gv_w_4 = _gv_w_4 + 1) begin : g_arb_data_in
													localparam w = _gv_w_4;
													// Trace: src/VX_scoreboard.sv:81:9
													assign arb_valid_in[w] = staging_if[w].valid && operands_ready[w];
													// Trace: src/VX_scoreboard.sv:82:9
													assign arb_data_in[w * 104+:104] = staging_if[w].data;
													// Trace: src/VX_scoreboard.sv:83:9
													assign staging_if[w].ready = arb_ready_in[w] && operands_ready[w];
												end
												// Trace: src/VX_scoreboard.sv:85:5
												VX_stream_arb #(
													.NUM_INPUTS(VX_gpu_pkg_PER_ISSUE_WARPS),
													.DATAW(DATAW),
													.ARBITER("C"),
													.OUT_BUF(3)
												) out_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(arb_valid_in),
													.ready_in(arb_ready_in),
													.data_in(arb_data_in),
													.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[105], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[102-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[98-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[67-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[65-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[61-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[24], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[23-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[17-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[11-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[5-:6]}),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.ready),
													.sel_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[104-:2])
												);
											end
											assign scoreboard.clk = clk;
											assign scoreboard.reset = reset;
											// Trace: src/VX_issue_slice.sv:31:5
											// expanded module instance: operands
											localparam _bbase_CD6E0_writeback_if = issue_id + _mbase_writeback_if;
											localparam _param_CD6E0_INSTANCE_ID = "";
											if (1) begin : operands
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_operands.sv:2:16
												localparam INSTANCE_ID = _param_CD6E0_INSTANCE_ID;
												// Trace: src/VX_operands.sv:3:15
												localparam NUM_BANKS = 4;
												// Trace: src/VX_operands.sv:4:15
												localparam OUT_BUF = 3;
												// Trace: src/VX_operands.sv:6:5
												wire clk;
												// Trace: src/VX_operands.sv:7:5
												wire reset;
												// Trace: src/VX_operands.sv:8:5
												localparam _mbase_writeback_if = _bbase_CD6E0_writeback_if;
												// Trace: src/VX_operands.sv:9:5
												// removed modport instance scoreboard_if
												// Trace: src/VX_operands.sv:10:5
												// removed modport instance operands_if
												// Trace: src/VX_operands.sv:12:5
												localparam NUM_SRC_OPDS = 3;
												// Trace: src/VX_operands.sv:13:5
												localparam REQ_SEL_BITS = 2;
												// Trace: src/VX_operands.sv:14:5
												localparam REQ_SEL_WIDTH = REQ_SEL_BITS;
												// Trace: src/VX_operands.sv:15:5
												localparam BANK_SEL_BITS = 2;
												// Trace: src/VX_operands.sv:16:5
												localparam BANK_SEL_WIDTH = BANK_SEL_BITS;
												// Trace: src/VX_operands.sv:17:5
												localparam PER_BANK_REGS = 16;
												// Trace: src/VX_operands.sv:18:5
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam VX_gpu_pkg_ISSUE_WIS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
												// removed localparam type VX_gpu_pkg_alu_args_t
												// removed localparam type VX_gpu_pkg_csr_args_t
												// removed localparam type VX_gpu_pkg_fpu_args_t
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam META_DATAW = 88;
												// Trace: src/VX_operands.sv:19:5
												localparam REGS_DATAW = 128;
												// Trace: src/VX_operands.sv:20:5
												localparam DATAW = 472;
												// Trace: src/VX_operands.sv:21:5
												localparam RAM_ADDRW = 8;
												// Trace: src/VX_operands.sv:22:5
												localparam PER_BANK_ADDRW = 6;
												// Trace: src/VX_operands.sv:23:5
												localparam XLEN_SIZE = 4;
												// Trace: src/VX_operands.sv:24:5
												localparam BYTEENW = 16;
												// Trace: src/VX_operands.sv:25:5
												wire [2:0] src_valid;
												// Trace: src/VX_operands.sv:26:5
												wire [2:0] req_valid_in;
												wire [2:0] req_ready_in;
												// Trace: src/VX_operands.sv:27:5
												wire [17:0] req_data_in;
												// Trace: src/VX_operands.sv:28:5
												wire [5:0] req_bank_idx;
												// Trace: src/VX_operands.sv:29:5
												wire [3:0] gpr_rd_valid;
												wire [3:0] gpr_rd_ready;
												// Trace: src/VX_operands.sv:30:5
												wire [3:0] gpr_rd_valid_st1;
												wire [3:0] gpr_rd_valid_st2;
												// Trace: src/VX_operands.sv:31:5
												wire [23:0] gpr_rd_addr;
												wire [23:0] gpr_rd_addr_st1;
												// Trace: src/VX_operands.sv:32:5
												wire [511:0] gpr_rd_data_st2;
												// Trace: src/VX_operands.sv:33:5
												wire [7:0] gpr_rd_req_idx;
												wire [7:0] gpr_rd_req_idx_st1;
												wire [7:0] gpr_rd_req_idx_st2;
												// Trace: src/VX_operands.sv:34:5
												wire pipe_ready_in;
												// Trace: src/VX_operands.sv:35:5
												wire pipe_valid_st1;
												wire pipe_ready_st1;
												// Trace: src/VX_operands.sv:36:5
												wire pipe_valid_st2;
												wire pipe_ready_st2;
												// Trace: src/VX_operands.sv:37:5
												wire [87:0] pipe_data;
												wire [87:0] pipe_data_st1;
												wire [87:0] pipe_data_st2;
												// Trace: src/VX_operands.sv:38:5
												reg [383:0] src_data_st2;
												reg [383:0] src_data_m_st2;
												// Trace: src/VX_operands.sv:39:5
												reg [2:0] data_fetched_st1;
												// Trace: src/VX_operands.sv:40:5
												reg has_collision_n;
												// Trace: src/VX_operands.sv:41:5
												wire has_collision_st1;
												// Trace: src/VX_operands.sv:42:5
												wire [17:0] src_opds;
												// Trace: src/VX_operands.sv:43:5
												assign src_opds = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[5-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[11-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[17-:6]};
												// Trace: src/VX_operands.sv:44:5
												genvar _gv_i_214;
												for (_gv_i_214 = 0; _gv_i_214 < NUM_SRC_OPDS; _gv_i_214 = _gv_i_214 + 1) begin : g_req_data_in
													localparam i = _gv_i_214;
													if (1) begin : g_wis
														// Trace: src/VX_operands.sv:46:13
														assign req_data_in[i * 6+:6] = {src_opds[(i * 6) + 5-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[104-:2]};
													end
												end
												// Trace: src/VX_operands.sv:51:5
												genvar _gv_i_215;
												for (_gv_i_215 = 0; _gv_i_215 < NUM_SRC_OPDS; _gv_i_215 = _gv_i_215 + 1) begin : g_req_bank_idx
													localparam i = _gv_i_215;
													if (1) begin : g_multibanks
														// Trace: src/VX_operands.sv:53:13
														assign req_bank_idx[i * 2+:2] = src_opds[(i * 6) + 1-:2];
													end
												end
												// Trace: src/VX_operands.sv:58:5
												genvar _gv_i_216;
												for (_gv_i_216 = 0; _gv_i_216 < NUM_SRC_OPDS; _gv_i_216 = _gv_i_216 + 1) begin : g_src_valid
													localparam i = _gv_i_216;
													// Trace: src/VX_operands.sv:59:9
													assign src_valid[i] = (src_opds[i * 6+:6] != 0) && ~data_fetched_st1[i];
												end
												// Trace: src/VX_operands.sv:61:5
												assign req_valid_in = {NUM_SRC_OPDS {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.valid}} & src_valid;
												// Trace: src/VX_operands.sv:62:5
												VX_stream_xbar #(
													.NUM_INPUTS(NUM_SRC_OPDS),
													.NUM_OUTPUTS(NUM_BANKS),
													.DATAW(PER_BANK_ADDRW),
													.ARBITER("P"),
													.PERF_CTR_BITS(44),
													.OUT_BUF(0)
												) req_xbar(
													.clk(clk),
													.reset(reset),
													.collisions(),
													.valid_in(req_valid_in),
													.data_in(req_data_in),
													.sel_in(req_bank_idx),
													.ready_in(req_ready_in),
													.valid_out(gpr_rd_valid),
													.data_out(gpr_rd_addr),
													.sel_out(gpr_rd_req_idx),
													.ready_out(gpr_rd_ready)
												);
												// Trace: src/VX_operands.sv:82:5
												assign gpr_rd_ready = {NUM_BANKS {pipe_ready_in}};
												// Trace: src/VX_operands.sv:83:5
												always @(*) begin
													// Trace: src/VX_operands.sv:84:9
													has_collision_n = 0;
													// Trace: src/VX_operands.sv:85:9
													begin : sv2v_autoblock_6
														// Trace: src/VX_operands.sv:85:14
														integer i;
														// Trace: src/VX_operands.sv:85:14
														for (i = 0; i < NUM_SRC_OPDS; i = i + 1)
															begin
																// Trace: src/VX_operands.sv:86:13
																begin : sv2v_autoblock_7
																	// Trace: src/VX_operands.sv:86:18
																	integer j;
																	// Trace: src/VX_operands.sv:86:18
																	for (j = 1; j < (NUM_SRC_OPDS - i); j = j + 1)
																		begin
																			// Trace: src/VX_operands.sv:87:17
																			has_collision_n = has_collision_n | ((src_valid[i] && src_valid[j + i]) && (req_bank_idx[i * 2+:2] == req_bank_idx[(j + i) * 2+:2]));
																		end
																end
															end
													end
												end
												// Trace: src/VX_operands.sv:93:5
												wire [2:0] req_fire_in = req_valid_in & req_ready_in;
												// Trace: src/VX_operands.sv:94:5
												assign pipe_data = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[104-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[102-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[98-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[24], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[67-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[65-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[61-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[23-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[105]};
												// Trace: src/VX_operands.sv:105:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.ready = pipe_ready_in && ~has_collision_n;
												// Trace: src/VX_operands.sv:106:5
												wire pipe_fire_st1 = pipe_valid_st1 && pipe_ready_st1;
												// Trace: src/VX_operands.sv:107:5
												wire pipe_fire_st2 = pipe_valid_st2 && pipe_ready_st2;
												// Trace: src/VX_operands.sv:108:5
												VX_pipe_buffer #(.DATAW(125)) pipe_reg1(
													.clk(clk),
													.reset(reset),
													.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.valid),
													.ready_in(pipe_ready_in),
													.data_in({gpr_rd_valid, pipe_data, has_collision_n, gpr_rd_addr, gpr_rd_req_idx}),
													.data_out({gpr_rd_valid_st1, pipe_data_st1, has_collision_st1, gpr_rd_addr_st1, gpr_rd_req_idx_st1}),
													.valid_out(pipe_valid_st1),
													.ready_out(pipe_ready_st1)
												);
												// Trace: src/VX_operands.sv:120:5
												always @(posedge clk)
													// Trace: src/VX_operands.sv:121:9
													if (reset || Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.ready)
														// Trace: src/VX_operands.sv:122:13
														data_fetched_st1 <= 0;
													else
														// Trace: src/VX_operands.sv:124:13
														data_fetched_st1 <= data_fetched_st1 | req_fire_in;
												// Trace: src/VX_operands.sv:127:5
												wire pipe_valid2_st1 = pipe_valid_st1 && ~has_collision_st1;
												// Trace: src/VX_operands.sv:128:5
												VX_pipe_buffer #(.DATAW(100)) pipe_reg2(
													.clk(clk),
													.reset(reset),
													.valid_in(pipe_valid2_st1),
													.ready_in(pipe_ready_st1),
													.data_in({gpr_rd_valid_st1, gpr_rd_req_idx_st1, pipe_data_st1}),
													.data_out({gpr_rd_valid_st2, gpr_rd_req_idx_st2, pipe_data_st2}),
													.valid_out(pipe_valid_st2),
													.ready_out(pipe_ready_st2)
												);
												// Trace: src/VX_operands.sv:140:5
												always @(*) begin
													// Trace: src/VX_operands.sv:141:9
													src_data_m_st2 = src_data_st2;
													// Trace: src/VX_operands.sv:142:9
													begin : sv2v_autoblock_8
														// Trace: src/VX_operands.sv:142:14
														integer b;
														// Trace: src/VX_operands.sv:142:14
														for (b = 0; b < NUM_BANKS; b = b + 1)
															begin
																// Trace: src/VX_operands.sv:143:13
																if (gpr_rd_valid_st2[b])
																	// Trace: src/VX_operands.sv:144:17
																	src_data_m_st2[gpr_rd_req_idx_st2[b * 2+:2] * 128+:128] = gpr_rd_data_st2[32 * (b * 4)+:128];
															end
													end
												end
												// Trace: src/VX_operands.sv:148:5
												always @(posedge clk)
													// Trace: src/VX_operands.sv:149:9
													if (reset || pipe_fire_st2)
														// Trace: src/VX_operands.sv:150:13
														src_data_st2 <= 0;
													else
														// Trace: src/VX_operands.sv:152:13
														src_data_st2 <= src_data_m_st2;
												// Trace: src/VX_operands.sv:155:5
												VX_elastic_buffer #(
													.DATAW(DATAW),
													.SIZE(2),
													.OUT_REG(1)
												) out_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(pipe_valid_st2),
													.ready_in(pipe_ready_st2),
													.data_in({pipe_data_st2, src_data_m_st2}),
													.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[470-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[468-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[464-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[390], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[433-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[431-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[427-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[389-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[471], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[127-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[255-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[383-:128]}),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.ready)
												);
												// Trace: src/VX_operands.sv:182:5
												wire [5:0] gpr_wr_addr;
												// Trace: src/VX_operands.sv:183:5
												if (1) begin : g_gpr_wr_addr
													// Trace: src/VX_operands.sv:184:9
													assign gpr_wr_addr = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[135:132], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[172-:2]};
												end
												// Trace: src/VX_operands.sv:188:5
												wire [1:0] gpr_wr_bank_idx;
												// Trace: src/VX_operands.sv:189:5
												if (1) begin : g_gpr_wr_bank_idx
													// Trace: src/VX_operands.sv:190:9
													assign gpr_wr_bank_idx = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[131:130];
												end
												// Trace: src/VX_operands.sv:194:5
												genvar _gv_b_1;
												for (_gv_b_1 = 0; _gv_b_1 < NUM_BANKS; _gv_b_1 = _gv_b_1 + 1) begin : g_gpr_rams
													localparam b = _gv_b_1;
													// Trace: src/VX_operands.sv:195:9
													wire gpr_wr_enabled;
													if (1) begin : g_gpr_wr_enabled_multibanks
														// Trace: src/VX_operands.sv:197:13
														assign gpr_wr_enabled = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].valid && (gpr_wr_bank_idx == sv2v_cast_2_signed(b));
													end
													// Trace: src/VX_operands.sv:202:9
													wire [15:0] wren;
													genvar _gv_i_217;
													for (_gv_i_217 = 0; _gv_i_217 < 4; _gv_i_217 = _gv_i_217 + 1) begin : g_wren
														localparam i = _gv_i_217;
														// Trace: src/VX_operands.sv:204:13
														assign wren[i * XLEN_SIZE+:XLEN_SIZE] = {XLEN_SIZE {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[167 + i]}};
													end
													// Trace: src/VX_operands.sv:206:9
													VX_dp_ram #(
														.DATAW(REGS_DATAW),
														.SIZE(64),
														.WRENW(BYTEENW),
														.OUT_REG(1),
														.RDW_MODE("U")
													) gpr_ram(
														.clk(clk),
														.reset(reset),
														.read(pipe_fire_st1),
														.wren(wren),
														.write(gpr_wr_enabled),
														.waddr(gpr_wr_addr),
														.wdata(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[129-:128]),
														.raddr(gpr_rd_addr_st1[b * 6+:6]),
														.rdata(gpr_rd_data_st2[32 * (b * 4)+:128])
													);
												end
											end
											assign operands.clk = clk;
											assign operands.reset = reset;
											// Trace: src/VX_issue_slice.sv:40:5
											// expanded module instance: dispatch
											localparam _bbase_1A128_dispatch_if = 0;
											localparam _param_1A128_INSTANCE_ID = "";
											if (1) begin : dispatch
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_dispatch.sv:2:16
												localparam INSTANCE_ID = _param_1A128_INSTANCE_ID;
												// Trace: src/VX_dispatch.sv:4:5
												wire clk;
												// Trace: src/VX_dispatch.sv:5:5
												wire reset;
												// Trace: src/VX_dispatch.sv:6:5
												// removed modport instance operands_if
												// Trace: src/VX_dispatch.sv:7:5
												localparam _mbase_dispatch_if = 0;
												// Trace: src/VX_dispatch.sv:9:5
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam VX_gpu_pkg_ISSUE_WIS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
												// removed localparam type VX_gpu_pkg_alu_args_t
												// removed localparam type VX_gpu_pkg_csr_args_t
												// removed localparam type VX_gpu_pkg_fpu_args_t
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam DATAW = 472;
												// Trace: src/VX_dispatch.sv:10:5
												wire [7:0] tids;
												// Trace: src/VX_dispatch.sv:11:5
												genvar _gv_i_151;
												for (_gv_i_151 = 0; _gv_i_151 < 4; _gv_i_151 = _gv_i_151 + 1) begin : g_tids
													localparam i = _gv_i_151;
													// Trace: src/VX_dispatch.sv:12:9
													assign tids[i * 2+:2] = sv2v_cast_2_signed(i);
												end
												// Trace: src/VX_dispatch.sv:14:5
												wire [1:0] last_active_tid;
												// Trace: src/VX_dispatch.sv:15:5
												VX_find_first #(
													.N(4),
													.DATAW(2),
													.REVERSE(1)
												) last_tid_select(
													.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[468-:4]),
													.data_in(tids),
													.data_out(last_active_tid),
													.valid_out()
												);
												// Trace: src/VX_dispatch.sv:25:5
												wire [3:0] operands_ready_in;
												// Trace: src/VX_dispatch.sv:26:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.ready = operands_ready_in[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[433-:2]];
												// Trace: src/VX_dispatch.sv:27:5
												genvar _gv_i_152;
												for (_gv_i_152 = 0; _gv_i_152 < 4; _gv_i_152 = _gv_i_152 + 1) begin : g_buffers
													localparam i = _gv_i_152;
													// Trace: src/VX_dispatch.sv:28:9
													VX_elastic_buffer #(
														.DATAW(DATAW),
														.SIZE(2),
														.OUT_REG(1)
													) buffer(
														.clk(clk),
														.reset(reset),
														.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.valid && (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[433-:2] == sv2v_cast_2_signed(i))),
														.ready_in(operands_ready_in[i]),
														.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[471], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[470-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[468-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[464-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[431-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[427-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[390], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[389-:6], last_active_tid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[383-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[255-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[127-:128]}),
														.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_dispatch_if[i + _mbase_dispatch_if].data),
														.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_dispatch_if[i + _mbase_dispatch_if].valid),
														.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_dispatch_if[i + _mbase_dispatch_if].ready)
													);
												end
											end
											assign dispatch.clk = clk;
											assign dispatch.reset = reset;
										end
										assign issue_slice.clk = clk;
										assign issue_slice.reset = reset;
										genvar _gv_ex_id_1;
										for (_gv_ex_id_1 = 0; _gv_ex_id_1 < 4; _gv_ex_id_1 = _gv_ex_id_1 + 1) begin : g_dispatch_if
											localparam ex_id = _gv_ex_id_1;
											// Trace: src/VX_issue.sv:45:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[((ex_id * 1) + issue_id) + _mbase_dispatch_if].valid = per_issue_dispatch_if[ex_id].valid;
											// Trace: src/VX_issue.sv:46:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[((ex_id * 1) + issue_id) + _mbase_dispatch_if].data = per_issue_dispatch_if[ex_id].data;
											// Trace: src/VX_issue.sv:47:5
											assign per_issue_dispatch_if[ex_id].ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[((ex_id * 1) + issue_id) + _mbase_dispatch_if].ready;
										end
									end
								end
								assign issue.clk = clk;
								assign issue.reset = reset;
								// Trace: src/VX_core.sv:79:5
								// expanded module instance: execute
								localparam _bbase_B78CA_lsu_mem_if = 0;
								localparam _bbase_B78CA_dispatch_if = 0;
								localparam _bbase_B78CA_commit_if = 0;
								localparam _bbase_B78CA_branch_ctl_if = 0;
								localparam _param_B78CA_INSTANCE_ID = "";
								localparam _param_B78CA_CORE_ID = CORE_ID;
								if (1) begin : execute
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_execute.sv:2:16
									localparam INSTANCE_ID = _param_B78CA_INSTANCE_ID;
									// Trace: src/VX_execute.sv:3:15
									localparam CORE_ID = _param_B78CA_CORE_ID;
									// Trace: src/VX_execute.sv:5:5
									wire clk;
									// Trace: src/VX_execute.sv:6:5
									wire reset;
									// Trace: src/VX_execute.sv:7:5
									// removed localparam type VX_gpu_pkg_base_dcrs_t
									wire [71:0] base_dcrs;
									// Trace: src/VX_execute.sv:8:5
									localparam _mbase_lsu_mem_if = 0;
									// Trace: src/VX_execute.sv:9:5
									localparam _mbase_dispatch_if = 0;
									// Trace: src/VX_execute.sv:10:5
									localparam _mbase_commit_if = 0;
									// Trace: src/VX_execute.sv:11:5
									// removed modport instance sched_csr_if
									// Trace: src/VX_execute.sv:12:5
									localparam _mbase_branch_ctl_if = 0;
									// Trace: src/VX_execute.sv:13:5
									// removed modport instance warp_ctl_if
									// Trace: src/VX_execute.sv:14:5
									// removed modport instance commit_csr_if
									// Trace: src/VX_execute.sv:16:5
									// expanded interface instance: fpu_csr_if
									genvar _arr_82930;
									for (_arr_82930 = 0; _arr_82930 <= 0; _arr_82930 = _arr_82930 + 1) begin : fpu_csr_if
										// removed import VX_fpu_pkg::*;
										// Trace: src/VX_fpu_csr_if.sv:2:5
										wire write_enable;
										// Trace: src/VX_fpu_csr_if.sv:3:5
										wire [1:0] write_wid;
										// Trace: src/VX_fpu_csr_if.sv:4:5
										// removed localparam type VX_fpu_pkg_fflags_t
										wire [4:0] write_fflags;
										// Trace: src/VX_fpu_csr_if.sv:5:5
										wire [1:0] read_wid;
										// Trace: src/VX_fpu_csr_if.sv:6:5
										wire [2:0] read_frm;
										// Trace: src/VX_fpu_csr_if.sv:7:5
										// Trace: src/VX_fpu_csr_if.sv:14:5
									end
									// Trace: src/VX_execute.sv:17:5
									// expanded module instance: alu_unit
									localparam _bbase_4B10A_dispatch_if = 0;
									localparam _bbase_4B10A_commit_if = 0;
									localparam _bbase_4B10A_branch_ctl_if = 0;
									localparam _param_4B10A_INSTANCE_ID = "";
									if (1) begin : alu_unit
										// Trace: src/VX_alu_unit.sv:2:16
										localparam INSTANCE_ID = _param_4B10A_INSTANCE_ID;
										// Trace: src/VX_alu_unit.sv:4:5
										wire clk;
										// Trace: src/VX_alu_unit.sv:5:5
										wire reset;
										// Trace: src/VX_alu_unit.sv:6:5
										localparam _mbase_dispatch_if = 0;
										// Trace: src/VX_alu_unit.sv:7:5
										localparam _mbase_commit_if = 0;
										// Trace: src/VX_alu_unit.sv:8:5
										localparam _mbase_branch_ctl_if = 0;
										// Trace: src/VX_alu_unit.sv:10:5
										localparam BLOCK_SIZE = 1;
										// Trace: src/VX_alu_unit.sv:11:5
										localparam NUM_LANES = 4;
										// Trace: src/VX_alu_unit.sv:12:5
										localparam PARTIAL_BW = 1'd0;
										// Trace: src/VX_alu_unit.sv:13:5
										localparam PE_COUNT = 2;
										// Trace: src/VX_alu_unit.sv:14:5
										localparam PE_SEL_BITS = 1;
										// Trace: src/VX_alu_unit.sv:15:5
										localparam PE_IDX_INT = 0;
										// Trace: src/VX_alu_unit.sv:16:5
										localparam PE_IDX_MDV = 1;
										// Trace: src/VX_alu_unit.sv:17:5
										// expanded interface instance: per_block_execute_if
										localparam _param_E2592_NUM_LANES = NUM_LANES;
										genvar _arr_E2592;
										for (_arr_E2592 = 0; _arr_E2592 <= 0; _arr_E2592 = _arr_E2592 + 1) begin : per_block_execute_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_execute_if.sv:2:15
											localparam NUM_LANES = _param_E2592_NUM_LANES;
											// Trace: src/VX_execute_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_execute_if.sv:5:5
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_execute_if.sv:22:5
											wire valid;
											// Trace: src/VX_execute_if.sv:23:5
											wire [474:0] data;
											// Trace: src/VX_execute_if.sv:24:5
											wire ready;
											// Trace: src/VX_execute_if.sv:25:5
											// Trace: src/VX_execute_if.sv:30:5
										end
										// Trace: src/VX_alu_unit.sv:20:5
										// expanded interface instance: per_block_commit_if
										localparam _param_98792_NUM_LANES = NUM_LANES;
										genvar _arr_98792;
										for (_arr_98792 = 0; _arr_98792 <= 0; _arr_98792 = _arr_98792 + 1) begin : per_block_commit_if
											// Trace: src/VX_commit_if.sv:2:15
											localparam NUM_LANES = _param_98792_NUM_LANES;
											// Trace: src/VX_commit_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_commit_if.sv:5:5
											// removed localparam type data_t
											// Trace: src/VX_commit_if.sv:17:5
											wire valid;
											// Trace: src/VX_commit_if.sv:18:5
											wire [175:0] data;
											// Trace: src/VX_commit_if.sv:19:5
											wire ready;
											// Trace: src/VX_commit_if.sv:20:5
											// Trace: src/VX_commit_if.sv:25:5
										end
										// Trace: src/VX_alu_unit.sv:23:5
										// expanded module instance: dispatch_unit
										localparam _bbase_2E16E_dispatch_if = 0;
										localparam _bbase_2E16E_execute_if = 0;
										localparam _param_2E16E_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_2E16E_NUM_LANES = NUM_LANES;
										localparam _param_2E16E_OUT_BUF = (PARTIAL_BW ? 3 : 0);
										if (1) begin : dispatch_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_dispatch_unit.sv:2:15
											localparam BLOCK_SIZE = _param_2E16E_BLOCK_SIZE;
											// Trace: src/VX_dispatch_unit.sv:3:15
											localparam NUM_LANES = _param_2E16E_NUM_LANES;
											// Trace: src/VX_dispatch_unit.sv:4:15
											localparam OUT_BUF = _param_2E16E_OUT_BUF;
											// Trace: src/VX_dispatch_unit.sv:5:15
											localparam MAX_FANOUT = 8;
											// Trace: src/VX_dispatch_unit.sv:7:5
											wire clk;
											// Trace: src/VX_dispatch_unit.sv:8:5
											wire reset;
											// Trace: src/VX_dispatch_unit.sv:9:5
											localparam _mbase_dispatch_if = 0;
											// Trace: src/VX_dispatch_unit.sv:10:5
											localparam _mbase_execute_if = 0;
											// Trace: src/VX_dispatch_unit.sv:12:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:13:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_dispatch_unit.sv:14:5
											localparam PID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:15:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:16:5
											localparam BATCH_COUNT = 1;
											// Trace: src/VX_dispatch_unit.sv:17:5
											localparam BATCH_COUNT_W = 1;
											// Trace: src/VX_dispatch_unit.sv:18:5
											localparam ISSUE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:19:5
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											localparam VX_gpu_pkg_ISSUE_WIS = 2;
											localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											localparam IN_DATAW = 472;
											// Trace: src/VX_dispatch_unit.sv:20:5
											localparam OUT_DATAW = 475;
											// Trace: src/VX_dispatch_unit.sv:21:5
											localparam FANOUT_ENABLE = 1'd0;
											// Trace: src/VX_dispatch_unit.sv:22:5
											localparam DATA_TMASK_OFF = 465;
											// Trace: src/VX_dispatch_unit.sv:23:5
											localparam DATA_REGS_OFF = 0;
											// Trace: src/VX_dispatch_unit.sv:24:5
											wire [0:0] dispatch_valid;
											// Trace: src/VX_dispatch_unit.sv:25:5
											wire [471:0] dispatch_data;
											// Trace: src/VX_dispatch_unit.sv:26:5
											wire [0:0] dispatch_ready;
											// Trace: src/VX_dispatch_unit.sv:27:5
											genvar _gv_i_96;
											for (_gv_i_96 = 0; _gv_i_96 < 1; _gv_i_96 = _gv_i_96 + 1) begin : g_dispatch_data
												localparam i = _gv_i_96;
												// Trace: src/VX_dispatch_unit.sv:28:9
												assign dispatch_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].valid;
												// Trace: src/VX_dispatch_unit.sv:29:9
												assign dispatch_data[i * 472+:472] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].data;
												// Trace: src/VX_dispatch_unit.sv:30:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].ready = dispatch_ready[i];
											end
											// Trace: src/VX_dispatch_unit.sv:32:5
											wire [0:0] block_ready;
											// Trace: src/VX_dispatch_unit.sv:33:5
											wire [3:0] block_tmask;
											// Trace: src/VX_dispatch_unit.sv:34:5
											wire [383:0] block_regs;
											// Trace: src/VX_dispatch_unit.sv:35:5
											wire [0:0] block_pid;
											// Trace: src/VX_dispatch_unit.sv:36:5
											wire [0:0] block_sop;
											// Trace: src/VX_dispatch_unit.sv:37:5
											wire [0:0] block_eop;
											// Trace: src/VX_dispatch_unit.sv:38:5
											wire [0:0] block_done;
											// Trace: src/VX_dispatch_unit.sv:39:5
											wire batch_done = &block_done;
											// Trace: src/VX_dispatch_unit.sv:40:5
											wire [0:0] batch_idx;
											// Trace: src/VX_dispatch_unit.sv:41:5
											if (1) begin : g_batch_idx_0
												// Trace: src/VX_dispatch_unit.sv:67:9
												assign batch_idx = 0;
											end
											// Trace: src/VX_dispatch_unit.sv:69:5
											wire [0:0] issue_indices;
											// Trace: src/VX_dispatch_unit.sv:70:5
											genvar _gv_block_idx_2;
											for (_gv_block_idx_2 = 0; _gv_block_idx_2 < BLOCK_SIZE; _gv_block_idx_2 = _gv_block_idx_2 + 1) begin : g_issue_indices
												localparam block_idx = _gv_block_idx_2;
												// Trace: src/VX_dispatch_unit.sv:71:9
												assign issue_indices[block_idx+:1] = sv2v_cast_1(batch_idx * BLOCK_SIZE) + sv2v_cast_1_signed(block_idx);
											end
											// Trace: src/VX_dispatch_unit.sv:73:5
											genvar _gv_block_idx_3;
											localparam VX_gpu_pkg_ISSUE_ISW = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											function [1:0] VX_gpu_pkg_wis_to_wid;
												// Trace: src/VX_gpu_pkg.sv:151:9
												input reg [1:0] wis;
												// Trace: src/VX_gpu_pkg.sv:152:9
												input reg [0:0] isw;
												// Trace: src/VX_gpu_pkg.sv:154:9
												begin
													// Trace: src/VX_gpu_pkg.sv:157:13
													VX_gpu_pkg_wis_to_wid = wis;
												end
											endfunction
											for (_gv_block_idx_3 = 0; _gv_block_idx_3 < BLOCK_SIZE; _gv_block_idx_3 = _gv_block_idx_3 + 1) begin : g_blocks
												localparam block_idx = _gv_block_idx_3;
												// Trace: src/VX_dispatch_unit.sv:74:9
												wire [0:0] issue_idx = issue_indices[block_idx+:1];
												// Trace: src/VX_dispatch_unit.sv:75:9
												wire valid_p;
												wire ready_p;
												if (1) begin : g_full_threads
													// Trace: src/VX_dispatch_unit.sv:168:13
													assign valid_p = dispatch_valid[issue_idx];
													// Trace: src/VX_dispatch_unit.sv:169:13
													assign block_tmask[block_idx * 4+:4] = dispatch_data[(issue_idx * 472) + DATA_TMASK_OFF+:4];
													// Trace: src/VX_dispatch_unit.sv:170:13
													assign block_regs[32 * ((block_idx * 3) * 4)+:128] = dispatch_data[(issue_idx * 472) + 256+:128];
													// Trace: src/VX_dispatch_unit.sv:171:13
													assign block_regs[32 * (((block_idx * 3) + 1) * 4)+:128] = dispatch_data[(issue_idx * 472) + 128+:128];
													// Trace: src/VX_dispatch_unit.sv:172:13
													assign block_regs[32 * (((block_idx * 3) + 2) * 4)+:128] = dispatch_data[issue_idx * 472+:128];
													// Trace: src/VX_dispatch_unit.sv:173:13
													assign block_pid[block_idx+:1] = 1'sb0;
													// Trace: src/VX_dispatch_unit.sv:174:13
													assign block_sop[block_idx] = 1'b1;
													// Trace: src/VX_dispatch_unit.sv:175:13
													assign block_eop[block_idx] = 1'b1;
													// Trace: src/VX_dispatch_unit.sv:176:13
													assign block_ready[block_idx] = ready_p;
													// Trace: src/VX_dispatch_unit.sv:177:13
													assign block_done[block_idx] = ready_p || ~valid_p;
												end
												// Trace: src/VX_dispatch_unit.sv:179:9
												wire [0:0] isw;
												if (1) begin : g_isw
													// Trace: src/VX_dispatch_unit.sv:187:13
													assign isw = block_idx;
												end
												// Trace: src/VX_dispatch_unit.sv:189:9
												wire [1:0] block_wid = VX_gpu_pkg_wis_to_wid(dispatch_data[(issue_idx * 472) + 469+:VX_gpu_pkg_ISSUE_WIS_W], isw);
												// Trace: src/VX_dispatch_unit.sv:190:9
												wire [474:0] execute_data;
												reg [474:0] execute_data_w;
												// Trace: src/VX_dispatch_unit.sv:191:9
												VX_elastic_buffer #(
													.DATAW(OUT_DATAW),
													.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
													.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
												) buf_out(
													.clk(clk),
													.reset(reset),
													.valid_in(valid_p),
													.ready_in(ready_p),
													.data_in({dispatch_data[(issue_idx * 472) + 471-:1], block_wid, block_tmask[block_idx * 4+:4], dispatch_data[(issue_idx * 472) + 464-:81], block_regs[32 * ((block_idx * 3) * 4)+:128], block_regs[32 * (((block_idx * 3) + 1) * 4)+:128], block_regs[32 * (((block_idx * 3) + 2) * 4)+:128], block_pid[block_idx+:1], block_sop[block_idx], block_eop[block_idx]}),
													.data_out(execute_data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[block_idx + _mbase_execute_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[block_idx + _mbase_execute_if].ready)
												);
												if (1) begin : g_execute_data_w_full
													// Trace: src/VX_dispatch_unit.sv:218:13
													always @(*) begin
														// Trace: src/VX_dispatch_unit.sv:219:17
														execute_data_w = execute_data;
														// Trace: src/VX_dispatch_unit.sv:220:17
														execute_data_w[2:0] = 3'b011;
													end
												end
												// Trace: src/VX_dispatch_unit.sv:223:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[block_idx + _mbase_execute_if].data = execute_data_w;
											end
											// Trace: src/VX_dispatch_unit.sv:225:5
											reg [0:0] ready_in;
											// Trace: src/VX_dispatch_unit.sv:226:5
											always @(*) begin
												// Trace: src/VX_dispatch_unit.sv:227:9
												ready_in = 0;
												// Trace: src/VX_dispatch_unit.sv:228:9
												begin : sv2v_autoblock_9
													// Trace: src/VX_dispatch_unit.sv:228:14
													integer block_idx;
													// Trace: src/VX_dispatch_unit.sv:228:14
													for (block_idx = 0; block_idx < BLOCK_SIZE; block_idx = block_idx + 1)
														begin
															// Trace: src/VX_dispatch_unit.sv:229:13
															ready_in[issue_indices[block_idx+:1]] = block_ready[block_idx] && block_eop[block_idx];
														end
												end
											end
											// Trace: src/VX_dispatch_unit.sv:232:5
											assign dispatch_ready = ready_in;
										end
										assign dispatch_unit.clk = clk;
										assign dispatch_unit.reset = reset;
										// Trace: src/VX_alu_unit.sv:33:5
										genvar _gv_block_idx_5;
										for (_gv_block_idx_5 = 0; _gv_block_idx_5 < BLOCK_SIZE; _gv_block_idx_5 = _gv_block_idx_5 + 1) begin : g_alus
											localparam block_idx = _gv_block_idx_5;
											// Trace: src/VX_alu_unit.sv:34:9
											// expanded interface instance: pe_execute_if
											localparam _param_C9035_NUM_LANES = NUM_LANES;
											genvar _arr_C9035;
											for (_arr_C9035 = 0; _arr_C9035 <= 1; _arr_C9035 = _arr_C9035 + 1) begin : pe_execute_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_execute_if.sv:2:15
												localparam NUM_LANES = _param_C9035_NUM_LANES;
												// Trace: src/VX_execute_if.sv:3:15
												localparam PID_WIDTH = 1;
												// Trace: src/VX_execute_if.sv:5:5
												// removed localparam type VX_gpu_pkg_alu_args_t
												// removed localparam type VX_gpu_pkg_csr_args_t
												// removed localparam type VX_gpu_pkg_fpu_args_t
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												// removed localparam type data_t
												// Trace: src/VX_execute_if.sv:22:5
												wire valid;
												// Trace: src/VX_execute_if.sv:23:5
												wire [474:0] data;
												// Trace: src/VX_execute_if.sv:24:5
												wire ready;
												// Trace: src/VX_execute_if.sv:25:5
												// Trace: src/VX_execute_if.sv:30:5
											end
											// Trace: src/VX_alu_unit.sv:37:9
											// expanded interface instance: pe_commit_if
											localparam _param_0FC39_NUM_LANES = NUM_LANES;
											genvar _arr_0FC39;
											for (_arr_0FC39 = 0; _arr_0FC39 <= 1; _arr_0FC39 = _arr_0FC39 + 1) begin : pe_commit_if
												// Trace: src/VX_commit_if.sv:2:15
												localparam NUM_LANES = _param_0FC39_NUM_LANES;
												// Trace: src/VX_commit_if.sv:3:15
												localparam PID_WIDTH = 1;
												// Trace: src/VX_commit_if.sv:5:5
												// removed localparam type data_t
												// Trace: src/VX_commit_if.sv:17:5
												wire valid;
												// Trace: src/VX_commit_if.sv:18:5
												wire [175:0] data;
												// Trace: src/VX_commit_if.sv:19:5
												wire ready;
												// Trace: src/VX_commit_if.sv:20:5
												// Trace: src/VX_commit_if.sv:25:5
											end
											// Trace: src/VX_alu_unit.sv:40:9
											reg [0:0] pe_select;
											// Trace: src/VX_alu_unit.sv:41:9
											always @(*) begin
												// Trace: src/VX_alu_unit.sv:42:13
												pe_select = PE_IDX_INT;
												// Trace: src/VX_alu_unit.sv:43:13
												if (per_block_execute_if[block_idx].data[429-:2] == 2)
													// Trace: src/VX_alu_unit.sv:44:17
													pe_select = PE_IDX_MDV;
											end
											// Trace: src/VX_alu_unit.sv:46:9
											// expanded module instance: pe_switch
											localparam _bbase_3D12E_execute_in_if = block_idx;
											localparam _bbase_3D12E_commit_out_if = block_idx;
											localparam _bbase_3D12E_execute_out_if = 0;
											localparam _bbase_3D12E_commit_in_if = 0;
											localparam _param_3D12E_PE_COUNT = PE_COUNT;
											localparam _param_3D12E_NUM_LANES = NUM_LANES;
											localparam _param_3D12E_ARBITER = "R";
											localparam _param_3D12E_REQ_OUT_BUF = 0;
											localparam _param_3D12E_RSP_OUT_BUF = (PARTIAL_BW ? 1 : 3);
											if (1) begin : pe_switch
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_pe_switch.sv:2:15
												localparam PE_COUNT = _param_3D12E_PE_COUNT;
												// Trace: src/VX_pe_switch.sv:3:15
												localparam NUM_LANES = _param_3D12E_NUM_LANES;
												// Trace: src/VX_pe_switch.sv:4:15
												localparam REQ_OUT_BUF = _param_3D12E_REQ_OUT_BUF;
												// Trace: src/VX_pe_switch.sv:5:15
												localparam RSP_OUT_BUF = _param_3D12E_RSP_OUT_BUF;
												// Trace: src/VX_pe_switch.sv:6:16
												localparam ARBITER = _param_3D12E_ARBITER;
												// Trace: src/VX_pe_switch.sv:7:15
												localparam PE_SEL_BITS = 1;
												// Trace: src/VX_pe_switch.sv:9:5
												wire clk;
												// Trace: src/VX_pe_switch.sv:10:5
												wire reset;
												// Trace: src/VX_pe_switch.sv:11:5
												wire [0:0] pe_sel;
												// Trace: src/VX_pe_switch.sv:12:5
												localparam _mbase_execute_in_if = _bbase_3D12E_execute_in_if;
												// Trace: src/VX_pe_switch.sv:13:5
												localparam _mbase_commit_out_if = _bbase_3D12E_commit_out_if;
												// Trace: src/VX_pe_switch.sv:14:5
												localparam _mbase_execute_out_if = 0;
												// Trace: src/VX_pe_switch.sv:15:5
												localparam _mbase_commit_in_if = 0;
												// Trace: src/VX_pe_switch.sv:17:5
												localparam PID_BITS = 0;
												// Trace: src/VX_pe_switch.sv:18:5
												localparam PID_WIDTH = 1;
												// Trace: src/VX_pe_switch.sv:19:5
												// removed localparam type VX_gpu_pkg_alu_args_t
												// removed localparam type VX_gpu_pkg_csr_args_t
												// removed localparam type VX_gpu_pkg_fpu_args_t
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam REQ_DATAW = 475;
												// Trace: src/VX_pe_switch.sv:20:5
												localparam RSP_DATAW = 176;
												// Trace: src/VX_pe_switch.sv:21:5
												wire [1:0] pe_req_valid;
												// Trace: src/VX_pe_switch.sv:22:5
												wire [949:0] pe_req_data;
												// Trace: src/VX_pe_switch.sv:23:5
												wire [1:0] pe_req_ready;
												// Trace: src/VX_pe_switch.sv:24:5
												VX_stream_switch #(
													.DATAW(REQ_DATAW),
													.NUM_INPUTS(1),
													.NUM_OUTPUTS(PE_COUNT),
													.OUT_BUF(REQ_OUT_BUF)
												) req_switch(
													.clk(clk),
													.reset(reset),
													.sel_in(pe_sel),
													.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[_mbase_execute_in_if].valid),
													.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[_mbase_execute_in_if].ready),
													.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[_mbase_execute_in_if].data),
													.data_out(pe_req_data),
													.valid_out(pe_req_valid),
													.ready_out(pe_req_ready)
												);
												// Trace: src/VX_pe_switch.sv:40:5
												genvar _gv_i_14;
												for (_gv_i_14 = 0; _gv_i_14 < PE_COUNT; _gv_i_14 = _gv_i_14 + 1) begin : g_execute_out_if
													localparam i = _gv_i_14;
													// Trace: src/VX_pe_switch.sv:41:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[i + _mbase_execute_out_if].valid = pe_req_valid[i];
													// Trace: src/VX_pe_switch.sv:42:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[i + _mbase_execute_out_if].data = pe_req_data[i * 475+:475];
													// Trace: src/VX_pe_switch.sv:43:9
													assign pe_req_ready[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[i + _mbase_execute_out_if].ready;
												end
												// Trace: src/VX_pe_switch.sv:45:5
												wire [1:0] pe_rsp_valid;
												// Trace: src/VX_pe_switch.sv:46:5
												wire [351:0] pe_rsp_data;
												// Trace: src/VX_pe_switch.sv:47:5
												wire [1:0] pe_rsp_ready;
												// Trace: src/VX_pe_switch.sv:48:5
												genvar _gv_i_15;
												for (_gv_i_15 = 0; _gv_i_15 < PE_COUNT; _gv_i_15 = _gv_i_15 + 1) begin : g_commit_in_if
													localparam i = _gv_i_15;
													// Trace: src/VX_pe_switch.sv:49:9
													assign pe_rsp_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[i + _mbase_commit_in_if].valid;
													// Trace: src/VX_pe_switch.sv:50:9
													assign pe_rsp_data[i * 176+:176] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[i + _mbase_commit_in_if].data;
													// Trace: src/VX_pe_switch.sv:51:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[i + _mbase_commit_in_if].ready = pe_rsp_ready[i];
												end
												// Trace: src/VX_pe_switch.sv:53:5
												VX_stream_arb #(
													.NUM_INPUTS(PE_COUNT),
													.DATAW(RSP_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(RSP_OUT_BUF)
												) rsp_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(pe_rsp_valid),
													.ready_in(pe_rsp_ready),
													.data_in(pe_rsp_data),
													.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_commit_if[_mbase_commit_out_if].data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_commit_if[_mbase_commit_out_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_commit_if[_mbase_commit_out_if].ready),
													.sel_out()
												);
											end
											assign pe_switch.clk = clk;
											assign pe_switch.reset = reset;
											assign pe_switch.pe_sel = pe_select;
											// Trace: src/VX_alu_unit.sv:61:9
											// expanded module instance: alu_int
											localparam _bbase_EF6D6_execute_if = PE_IDX_INT;
											localparam _bbase_EF6D6_branch_ctl_if = block_idx + _mbase_branch_ctl_if;
											localparam _bbase_EF6D6_commit_if = PE_IDX_INT;
											localparam _param_EF6D6_INSTANCE_ID = "";
											localparam _param_EF6D6_BLOCK_IDX = block_idx;
											localparam _param_EF6D6_NUM_LANES = NUM_LANES;
											if (1) begin : alu_int
												// Trace: src/VX_alu_int.sv:2:16
												localparam INSTANCE_ID = _param_EF6D6_INSTANCE_ID;
												// Trace: src/VX_alu_int.sv:3:15
												localparam BLOCK_IDX = _param_EF6D6_BLOCK_IDX;
												// Trace: src/VX_alu_int.sv:4:15
												localparam NUM_LANES = _param_EF6D6_NUM_LANES;
												// Trace: src/VX_alu_int.sv:6:5
												wire clk;
												// Trace: src/VX_alu_int.sv:7:5
												wire reset;
												// Trace: src/VX_alu_int.sv:8:5
												localparam _mbase_execute_if = _bbase_EF6D6_execute_if;
												// Trace: src/VX_alu_int.sv:9:5
												localparam _mbase_commit_if = _bbase_EF6D6_commit_if;
												// Trace: src/VX_alu_int.sv:10:5
												localparam _mbase_branch_ctl_if = _bbase_EF6D6_branch_ctl_if;
												// Trace: src/VX_alu_int.sv:12:5
												localparam LANE_BITS = 2;
												// Trace: src/VX_alu_int.sv:13:5
												localparam LANE_WIDTH = LANE_BITS;
												// Trace: src/VX_alu_int.sv:14:5
												localparam PID_BITS = 0;
												// Trace: src/VX_alu_int.sv:15:5
												localparam PID_WIDTH = 1;
												// Trace: src/VX_alu_int.sv:16:5
												localparam SHIFT_IMM_BITS = 5;
												// Trace: src/VX_alu_int.sv:17:5
												wire [127:0] add_result;
												// Trace: src/VX_alu_int.sv:18:5
												wire [131:0] sub_result;
												// Trace: src/VX_alu_int.sv:19:5
												reg [127:0] shr_zic_result;
												// Trace: src/VX_alu_int.sv:20:5
												reg [127:0] msc_result;
												// Trace: src/VX_alu_int.sv:21:5
												wire [127:0] add_result_w;
												// Trace: src/VX_alu_int.sv:22:5
												wire [127:0] sub_result_w;
												// Trace: src/VX_alu_int.sv:23:5
												wire [127:0] shr_result_w;
												// Trace: src/VX_alu_int.sv:24:5
												reg [127:0] msc_result_w;
												// Trace: src/VX_alu_int.sv:25:5
												reg [127:0] alu_result;
												// Trace: src/VX_alu_int.sv:26:5
												wire [127:0] alu_result_r;
												// Trace: src/VX_alu_int.sv:27:5
												wire is_alu_w = 0;
												// Trace: src/VX_alu_int.sv:28:5
												wire [3:0] alu_op = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[436-:4];
												// Trace: src/VX_alu_int.sv:29:5
												wire [3:0] br_op = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[436-:4];
												// Trace: src/VX_alu_int.sv:30:5
												wire is_br_op = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[429-:2] == 1;
												// Trace: src/VX_alu_int.sv:31:5
												wire is_sub_op = alu_op[1];
												// Trace: src/VX_alu_int.sv:32:5
												wire is_signed = alu_op[0];
												// Trace: src/VX_alu_int.sv:33:5
												wire [1:0] op_class = (is_br_op ? {1'b0, ~alu_op[3]} : alu_op[3:2]);
												// Trace: src/VX_alu_int.sv:34:5
												wire [127:0] alu_in1 = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[386-:128];
												// Trace: src/VX_alu_int.sv:35:5
												wire [127:0] alu_in2 = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[258-:128];
												// Trace: src/VX_alu_int.sv:36:5
												wire [127:0] alu_in1_PC = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[432] ? {NUM_LANES {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[467-:31], 1'd0}} : alu_in1);
												// Trace: src/VX_alu_int.sv:37:5
												wire [127:0] alu_in2_imm = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[431] ? {NUM_LANES {{Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[427], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[426:396]}}} : alu_in2);
												// Trace: src/VX_alu_int.sv:38:5
												wire [127:0] alu_in2_br = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[431] && ~is_br_op ? {NUM_LANES {{Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[427], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[426:396]}}} : alu_in2);
												// Trace: src/VX_alu_int.sv:39:5
												genvar _gv_i_8;
												for (_gv_i_8 = 0; _gv_i_8 < NUM_LANES; _gv_i_8 = _gv_i_8 + 1) begin : g_add_result
													localparam i = _gv_i_8;
													// Trace: src/VX_alu_int.sv:40:9
													assign add_result[i * 32+:32] = alu_in1_PC[i * 32+:32] + alu_in2_imm[i * 32+:32];
													// Trace: src/VX_alu_int.sv:41:9
													assign add_result_w[i * 32+:32] = sv2v_cast_32_signed($signed(alu_in1[(i * 32) + 31-:32] + alu_in2_imm[(i * 32) + 31-:32]));
												end
												// Trace: src/VX_alu_int.sv:43:5
												genvar _gv_i_9;
												for (_gv_i_9 = 0; _gv_i_9 < NUM_LANES; _gv_i_9 = _gv_i_9 + 1) begin : g_sub_result
													localparam i = _gv_i_9;
													// Trace: src/VX_alu_int.sv:44:9
													wire [32:0] sub_in1 = {is_signed & alu_in1[(i * 32) + 31], alu_in1[i * 32+:32]};
													// Trace: src/VX_alu_int.sv:45:9
													wire [32:0] sub_in2 = {is_signed & alu_in2_br[(i * 32) + 31], alu_in2_br[i * 32+:32]};
													// Trace: src/VX_alu_int.sv:46:9
													assign sub_result[i * 33+:33] = sub_in1 - sub_in2;
													// Trace: src/VX_alu_int.sv:47:9
													assign sub_result_w[i * 32+:32] = sv2v_cast_32_signed($signed(alu_in1[(i * 32) + 31-:32] - alu_in2_imm[(i * 32) + 31-:32]));
												end
												// Trace: src/VX_alu_int.sv:49:5
												genvar _gv_i_10;
												for (_gv_i_10 = 0; _gv_i_10 < NUM_LANES; _gv_i_10 = _gv_i_10 + 1) begin : g_shr_result
													localparam i = _gv_i_10;
													// Trace: src/VX_alu_int.sv:50:9
													wire [32:0] shr_in1 = {is_signed && alu_in1[(i * 32) + 31], alu_in1[i * 32+:32]};
													// Trace: src/VX_alu_int.sv:51:9
													always @(*)
														// Trace: src/VX_alu_int.sv:52:13
														case (alu_op[1:0])
															2'b10, 2'b11:
																// Trace: src/VX_alu_int.sv:54:21
																shr_zic_result[i * 32+:32] = alu_in1[i * 32+:32] & {32 {alu_op[0] ^ |alu_in2[i * 32+:32]}};
															default:
																// Trace: src/VX_alu_int.sv:57:21
																shr_zic_result[i * 32+:32] = sv2v_cast_32_signed($signed(shr_in1) >>> alu_in2_imm[(i * 32) + 4-:5]);
														endcase
													// Trace: src/VX_alu_int.sv:61:9
													wire [32:0] shr_in1_w = {is_signed && alu_in1[(i * 32) + 31], alu_in1[(i * 32) + 31-:32]};
													// Trace: src/VX_alu_int.sv:62:9
													wire [31:0] shr_res_w = sv2v_cast_32_signed($signed(shr_in1_w) >>> alu_in2_imm[(i * 32) + 4-:5]);
													// Trace: src/VX_alu_int.sv:63:9
													assign shr_result_w[i * 32+:32] = sv2v_cast_32_signed($signed(shr_res_w));
												end
												// Trace: src/VX_alu_int.sv:65:5
												genvar _gv_i_11;
												for (_gv_i_11 = 0; _gv_i_11 < NUM_LANES; _gv_i_11 = _gv_i_11 + 1) begin : g_msc_result
													localparam i = _gv_i_11;
													// Trace: src/VX_alu_int.sv:66:9
													always @(*)
														// Trace: src/VX_alu_int.sv:67:13
														case (alu_op[1:0])
															2'b00:
																// Trace: src/VX_alu_int.sv:68:24
																msc_result[i * 32+:32] = alu_in1[i * 32+:32] & alu_in2_imm[i * 32+:32];
															2'b01:
																// Trace: src/VX_alu_int.sv:69:24
																msc_result[i * 32+:32] = alu_in1[i * 32+:32] | alu_in2_imm[i * 32+:32];
															2'b10:
																// Trace: src/VX_alu_int.sv:70:24
																msc_result[i * 32+:32] = alu_in1[i * 32+:32] ^ alu_in2_imm[i * 32+:32];
															2'b11:
																// Trace: src/VX_alu_int.sv:71:24
																msc_result[i * 32+:32] = alu_in1[i * 32+:32] << alu_in2_imm[(i * 32) + 4-:5];
														endcase
													// Trace: src/VX_alu_int.sv:74:9
													wire [32:1] sv2v_tmp_4E506;
													assign sv2v_tmp_4E506 = sv2v_cast_32_signed($signed(alu_in1[(i * 32) + 31-:32] << alu_in2_imm[(i * 32) + 4-:5]));
													always @(*) msc_result_w[i * 32+:32] = sv2v_tmp_4E506;
												end
												// Trace: src/VX_alu_int.sv:76:5
												genvar _gv_i_12;
												for (_gv_i_12 = 0; _gv_i_12 < NUM_LANES; _gv_i_12 = _gv_i_12 + 1) begin : g_alu_result
													localparam i = _gv_i_12;
													// Trace: src/VX_alu_int.sv:77:9
													wire [31:0] slt_br_result = sv2v_cast_32({is_br_op && ~(|sub_result[(i * 33) + 31-:32]), sub_result[(i * 33) + 32]});
													// Trace: src/VX_alu_int.sv:78:9
													wire [31:0] sub_slt_br_result = (is_sub_op && ~is_br_op ? sub_result[(i * 33) + 31-:32] : slt_br_result);
													// Trace: src/VX_alu_int.sv:79:9
													always @(*)
														// Trace: src/VX_alu_int.sv:80:13
														case ({is_alu_w, op_class})
															3'b000:
																// Trace: src/VX_alu_int.sv:81:25
																alu_result[i * 32+:32] = add_result[i * 32+:32];
															3'b001:
																// Trace: src/VX_alu_int.sv:82:25
																alu_result[i * 32+:32] = sub_slt_br_result;
															3'b010:
																// Trace: src/VX_alu_int.sv:83:25
																alu_result[i * 32+:32] = shr_zic_result[i * 32+:32];
															3'b011:
																// Trace: src/VX_alu_int.sv:84:25
																alu_result[i * 32+:32] = msc_result[i * 32+:32];
															3'b100:
																// Trace: src/VX_alu_int.sv:85:25
																alu_result[i * 32+:32] = add_result_w[i * 32+:32];
															3'b101:
																// Trace: src/VX_alu_int.sv:86:25
																alu_result[i * 32+:32] = sub_result_w[i * 32+:32];
															3'b110:
																// Trace: src/VX_alu_int.sv:87:25
																alu_result[i * 32+:32] = shr_result_w[i * 32+:32];
															3'b111:
																// Trace: src/VX_alu_int.sv:88:25
																alu_result[i * 32+:32] = msc_result_w[i * 32+:32];
														endcase
												end
												// Trace: src/VX_alu_int.sv:92:5
												wire [30:0] PC_r;
												// Trace: src/VX_alu_int.sv:93:5
												wire [3:0] br_op_r;
												// Trace: src/VX_alu_int.sv:94:5
												wire [30:0] cbr_dest;
												wire [30:0] cbr_dest_r;
												// Trace: src/VX_alu_int.sv:95:5
												wire [1:0] tid;
												wire [1:0] tid_r;
												// Trace: src/VX_alu_int.sv:96:5
												wire is_br_op_r;
												// Trace: src/VX_alu_int.sv:97:5
												assign cbr_dest = add_result[1+:31];
												// Trace: src/VX_alu_int.sv:98:5
												if (1) begin : g_tid
													// Trace: src/VX_alu_int.sv:99:9
													assign tid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[387+:LANE_BITS];
												end
												// Trace: src/VX_alu_int.sv:103:5
												VX_elastic_buffer #(.DATAW(214)) rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].valid),
													.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].ready),
													.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[474], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[473-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[471-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[394-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[395], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[0], alu_result, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[467-:31], cbr_dest, is_br_op, br_op, tid}),
													.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[175], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[174-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[172-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[136-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[137], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[0], alu_result_r, PC_r, cbr_dest_r, is_br_op_r, br_op_r, tid_r}),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].ready)
												);
												// Trace: src/VX_alu_int.sv:115:5
												wire is_br_neg = br_op_r[1];
												// Trace: src/VX_alu_int.sv:116:5
												wire is_br_less = br_op_r[2];
												// Trace: src/VX_alu_int.sv:117:5
												wire is_br_static = br_op_r[3];
												// Trace: src/VX_alu_int.sv:118:5
												wire [31:0] br_result = alu_result_r[tid_r * 32+:32];
												// Trace: src/VX_alu_int.sv:119:5
												wire is_less = br_result[0];
												// Trace: src/VX_alu_int.sv:120:5
												wire is_equal = br_result[1];
												// Trace: src/VX_alu_int.sv:121:5
												wire br_enable = ((is_br_op_r && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].valid) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].ready) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[0];
												// Trace: src/VX_alu_int.sv:122:5
												wire br_taken = ((is_br_less ? is_less : is_equal) ^ is_br_neg) | is_br_static;
												// Trace: src/VX_alu_int.sv:123:5
												wire [30:0] br_dest = (is_br_static ? br_result[1+:31] : cbr_dest_r);
												// Trace: src/VX_alu_int.sv:124:5
												wire [1:0] br_wid;
												// Trace: src/VX_alu_int.sv:126:5
												if (1) begin : genblk7
													// Trace: src/VX_alu_int.sv:133:9
													assign br_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[174-:2];
												end
												// Trace: src/VX_alu_int.sv:136:5
												VX_pipe_register #(.DATAW(35)) branch_reg(
													.clk(clk),
													.reset(reset),
													.enable(1'b1),
													.data_in({br_enable, br_wid, br_taken, br_dest}),
													.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[_mbase_branch_ctl_if].valid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[_mbase_branch_ctl_if].wid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[_mbase_branch_ctl_if].taken, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[_mbase_branch_ctl_if].dest})
												);
												// Trace: src/VX_alu_int.sv:145:5
												genvar _gv_i_13;
												for (_gv_i_13 = 0; _gv_i_13 < NUM_LANES; _gv_i_13 = _gv_i_13 + 1) begin : g_commit
													localparam i = _gv_i_13;
													// Trace: src/VX_alu_int.sv:146:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[3 + (i * 32)+:32] = (is_br_op_r && is_br_static ? {PC_r + 31'sd2, 1'd0} : alu_result_r[i * 32+:32]);
												end
												// Trace: src/VX_alu_int.sv:148:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[168-:31] = PC_r;
											end
											assign alu_int.clk = clk;
											assign alu_int.reset = reset;
											// Trace: src/VX_alu_unit.sv:72:9
											// expanded module instance: muldiv_unit
											localparam _bbase_50917_execute_if = PE_IDX_MDV;
											localparam _bbase_50917_commit_if = PE_IDX_MDV;
											localparam _param_50917_INSTANCE_ID = "";
											localparam _param_50917_NUM_LANES = NUM_LANES;
											if (1) begin : muldiv_unit
												// Trace: src/VX_alu_muldiv.sv:2:16
												localparam INSTANCE_ID = _param_50917_INSTANCE_ID;
												// Trace: src/VX_alu_muldiv.sv:3:15
												localparam NUM_LANES = _param_50917_NUM_LANES;
												// Trace: src/VX_alu_muldiv.sv:5:5
												wire clk;
												// Trace: src/VX_alu_muldiv.sv:6:5
												wire reset;
												// Trace: src/VX_alu_muldiv.sv:7:5
												localparam _mbase_execute_if = _bbase_50917_execute_if;
												// Trace: src/VX_alu_muldiv.sv:8:5
												localparam _mbase_commit_if = _bbase_50917_commit_if;
												// Trace: src/VX_alu_muldiv.sv:10:5
												localparam PID_BITS = 0;
												// Trace: src/VX_alu_muldiv.sv:11:5
												localparam PID_WIDTH = 1;
												// Trace: src/VX_alu_muldiv.sv:12:5
												localparam TAG_WIDTH = 48;
												// Trace: src/VX_alu_muldiv.sv:13:5
												wire [2:0] muldiv_op = sv2v_cast_3(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[436-:4]);
												// Trace: src/VX_alu_muldiv.sv:14:5
												wire is_mulx_op = ~muldiv_op[2];
												// Trace: src/VX_alu_muldiv.sv:15:5
												wire is_signed_op = ~muldiv_op[0];
												// Trace: src/VX_alu_muldiv.sv:16:5
												wire is_alu_w = 0;
												// Trace: src/VX_alu_muldiv.sv:17:5
												wire [127:0] mul_result_out;
												// Trace: src/VX_alu_muldiv.sv:18:5
												wire [0:0] mul_uuid_out;
												// Trace: src/VX_alu_muldiv.sv:19:5
												wire [1:0] mul_wid_out;
												// Trace: src/VX_alu_muldiv.sv:20:5
												wire [3:0] mul_tmask_out;
												// Trace: src/VX_alu_muldiv.sv:21:5
												wire [30:0] mul_PC_out;
												// Trace: src/VX_alu_muldiv.sv:22:5
												wire [5:0] mul_rd_out;
												// Trace: src/VX_alu_muldiv.sv:23:5
												wire mul_wb_out;
												// Trace: src/VX_alu_muldiv.sv:24:5
												wire [0:0] mul_pid_out;
												// Trace: src/VX_alu_muldiv.sv:25:5
												wire mul_sop_out;
												wire mul_eop_out;
												// Trace: src/VX_alu_muldiv.sv:26:5
												wire mul_valid_in = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].valid && is_mulx_op;
												// Trace: src/VX_alu_muldiv.sv:27:5
												wire mul_ready_in;
												// Trace: src/VX_alu_muldiv.sv:28:5
												wire mul_valid_out;
												// Trace: src/VX_alu_muldiv.sv:29:5
												wire mul_ready_out;
												// Trace: src/VX_alu_muldiv.sv:30:5
												wire is_mulh_in = muldiv_op[1:0] != 0;
												// Trace: src/VX_alu_muldiv.sv:31:5
												wire is_signed_mul_a = muldiv_op[1:0] != 1;
												// Trace: src/VX_alu_muldiv.sv:32:5
												wire is_signed_mul_b = is_signed_op;
												// Trace: src/VX_alu_muldiv.sv:33:5
												wire [263:0] mul_result_tmp;
												// Trace: src/VX_alu_muldiv.sv:34:5
												wire is_mulh_out;
												// Trace: src/VX_alu_muldiv.sv:35:5
												wire is_mul_w_out;
												// Trace: src/VX_alu_muldiv.sv:36:5
												genvar _gv_i_186;
												for (_gv_i_186 = 0; _gv_i_186 < NUM_LANES; _gv_i_186 = _gv_i_186 + 1) begin : g_multiplier
													localparam i = _gv_i_186;
													// Trace: src/VX_alu_muldiv.sv:37:9
													wire [32:0] mul_in1 = {is_signed_mul_a && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[259 + ((i * 32) + 31)], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[259 + (i * 32)+:32]};
													// Trace: src/VX_alu_muldiv.sv:38:9
													wire [32:0] mul_in2 = {is_signed_mul_b && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[131 + ((i * 32) + 31)], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[131 + (i * 32)+:32]};
													// Trace: src/VX_alu_muldiv.sv:39:9
													VX_multiplier #(
														.A_WIDTH(33),
														.B_WIDTH(33),
														.R_WIDTH(66),
														.SIGNED(1),
														.LATENCY(4)
													) multiplier(
														.clk(clk),
														.enable(mul_ready_in),
														.dataa(mul_in1),
														.datab(mul_in2),
														.result(mul_result_tmp[i * 66+:66])
													);
												end
												// Trace: src/VX_alu_muldiv.sv:53:5
												VX_shift_register #(
													.DATAW(51),
													.DEPTH(4),
													.RESETW(1)
												) mul_shift_reg(
													.clk(clk),
													.reset(reset),
													.enable(mul_ready_in),
													.data_in({mul_valid_in, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[474], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[473-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[471-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[467-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[394-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[395], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[0], is_mulh_in, is_alu_w}),
													.data_out({mul_valid_out, mul_uuid_out, mul_wid_out, mul_tmask_out, mul_PC_out, mul_rd_out, mul_wb_out, mul_pid_out, mul_sop_out, mul_eop_out, is_mulh_out, is_mul_w_out})
												);
												// Trace: src/VX_alu_muldiv.sv:64:5
												assign mul_ready_in = mul_ready_out || ~mul_valid_out;
												// Trace: src/VX_alu_muldiv.sv:65:5
												genvar _gv_i_187;
												for (_gv_i_187 = 0; _gv_i_187 < NUM_LANES; _gv_i_187 = _gv_i_187 + 1) begin : g_mul_result_out
													localparam i = _gv_i_187;
													// Trace: src/VX_alu_muldiv.sv:66:9
													assign mul_result_out[i * 32+:32] = (is_mulh_out ? mul_result_tmp[(i * 66) + 63-:32] : mul_result_tmp[(i * 66) + 31-:32]);
												end
												// Trace: src/VX_alu_muldiv.sv:68:5
												wire [127:0] div_result_out;
												// Trace: src/VX_alu_muldiv.sv:69:5
												wire [0:0] div_uuid_out;
												// Trace: src/VX_alu_muldiv.sv:70:5
												wire [1:0] div_wid_out;
												// Trace: src/VX_alu_muldiv.sv:71:5
												wire [3:0] div_tmask_out;
												// Trace: src/VX_alu_muldiv.sv:72:5
												wire [30:0] div_PC_out;
												// Trace: src/VX_alu_muldiv.sv:73:5
												wire [5:0] div_rd_out;
												// Trace: src/VX_alu_muldiv.sv:74:5
												wire div_wb_out;
												// Trace: src/VX_alu_muldiv.sv:75:5
												wire [0:0] div_pid_out;
												// Trace: src/VX_alu_muldiv.sv:76:5
												wire div_sop_out;
												wire div_eop_out;
												// Trace: src/VX_alu_muldiv.sv:77:5
												wire is_rem_op = muldiv_op[1];
												// Trace: src/VX_alu_muldiv.sv:78:5
												wire div_valid_in = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].valid && ~is_mulx_op;
												// Trace: src/VX_alu_muldiv.sv:79:5
												wire div_ready_in;
												// Trace: src/VX_alu_muldiv.sv:80:5
												wire div_valid_out;
												// Trace: src/VX_alu_muldiv.sv:81:5
												wire div_ready_out;
												// Trace: src/VX_alu_muldiv.sv:82:5
												wire [127:0] div_in1;
												// Trace: src/VX_alu_muldiv.sv:83:5
												wire [127:0] div_in2;
												// Trace: src/VX_alu_muldiv.sv:84:5
												genvar _gv_i_188;
												for (_gv_i_188 = 0; _gv_i_188 < NUM_LANES; _gv_i_188 = _gv_i_188 + 1) begin : g_div_in
													localparam i = _gv_i_188;
													// Trace: src/VX_alu_muldiv.sv:85:9
													assign div_in1[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[259 + (i * 32)+:32];
													// Trace: src/VX_alu_muldiv.sv:86:9
													assign div_in2[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[131 + (i * 32)+:32];
												end
												// Trace: src/VX_alu_muldiv.sv:88:5
												wire [127:0] div_quotient;
												wire [127:0] div_remainder;
												// Trace: src/VX_alu_muldiv.sv:89:5
												wire is_rem_op_out;
												// Trace: src/VX_alu_muldiv.sv:90:5
												wire is_div_w_out;
												// Trace: src/VX_alu_muldiv.sv:91:5
												wire div_strode;
												// Trace: src/VX_alu_muldiv.sv:92:5
												wire div_busy;
												// Trace: src/VX_alu_muldiv.sv:93:5
												VX_elastic_adapter div_elastic_adapter(
													.clk(clk),
													.reset(reset),
													.valid_in(div_valid_in),
													.ready_in(div_ready_in),
													.valid_out(div_valid_out),
													.ready_out(div_ready_out),
													.strobe(div_strode),
													.busy(div_busy)
												);
												// Trace: src/VX_alu_muldiv.sv:103:5
												VX_serial_div #(
													.WIDTHN(32),
													.WIDTHD(32),
													.WIDTHQ(32),
													.WIDTHR(32),
													.LANES(NUM_LANES)
												) serial_div(
													.clk(clk),
													.reset(reset),
													.strobe(div_strode),
													.busy(div_busy),
													.is_signed(is_signed_op),
													.numer(div_in1),
													.denom(div_in2),
													.quotient(div_quotient),
													.remainder(div_remainder)
												);
												// Trace: src/VX_alu_muldiv.sv:120:5
												reg [49:0] div_tag_r;
												// Trace: src/VX_alu_muldiv.sv:121:5
												always @(posedge clk)
													// Trace: src/VX_alu_muldiv.sv:122:9
													if (div_valid_in && div_ready_in)
														// Trace: src/VX_alu_muldiv.sv:123:13
														div_tag_r <= {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[474], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[473-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[471-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[467-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[394-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[395], is_rem_op, is_alu_w, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].data[0]};
												// Trace: src/VX_alu_muldiv.sv:126:5
												assign {div_uuid_out, div_wid_out, div_tmask_out, div_PC_out, div_rd_out, div_wb_out, is_rem_op_out, is_div_w_out, div_pid_out, div_sop_out, div_eop_out} = div_tag_r;
												// Trace: src/VX_alu_muldiv.sv:127:5
												genvar _gv_i_189;
												for (_gv_i_189 = 0; _gv_i_189 < NUM_LANES; _gv_i_189 = _gv_i_189 + 1) begin : g_div_result_out
													localparam i = _gv_i_189;
													// Trace: src/VX_alu_muldiv.sv:128:9
													assign div_result_out[i * 32+:32] = (is_rem_op_out ? div_remainder[i * 32+:32] : div_quotient[i * 32+:32]);
												end
												// Trace: src/VX_alu_muldiv.sv:130:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_execute_if[_mbase_execute_if].ready = (is_mulx_op ? mul_ready_in : div_ready_in);
												// Trace: src/VX_alu_muldiv.sv:131:5
												VX_stream_arb #(
													.NUM_INPUTS(2),
													.DATAW(176),
													.ARBITER("P"),
													.OUT_BUF(2)
												) rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in({div_valid_out, mul_valid_out}),
													.ready_in({div_ready_out, mul_ready_out}),
													.data_in({div_uuid_out, div_wid_out, div_tmask_out, div_PC_out, div_rd_out, div_wb_out, div_pid_out, div_sop_out, div_eop_out, div_result_out, mul_uuid_out, mul_wid_out, mul_tmask_out, mul_PC_out, mul_rd_out, mul_wb_out, mul_pid_out, mul_sop_out, mul_eop_out, mul_result_out}),
													.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[175], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[174-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[172-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[168-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[136-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[137], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[0], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].data[130-:128]}),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_alus[_gv_block_idx_5].pe_commit_if[_mbase_commit_if].ready),
													.sel_out()
												);
											end
											assign muldiv_unit.clk = clk;
											assign muldiv_unit.reset = reset;
										end
										// Trace: src/VX_alu_unit.sv:82:5
										// expanded module instance: gather_unit
										localparam _bbase_8E516_commit_in_if = 0;
										localparam _bbase_8E516_commit_out_if = 0;
										localparam _param_8E516_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_8E516_NUM_LANES = NUM_LANES;
										localparam _param_8E516_OUT_BUF = (PARTIAL_BW ? 3 : 0);
										if (1) begin : gather_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_gather_unit.sv:2:15
											localparam BLOCK_SIZE = _param_8E516_BLOCK_SIZE;
											// Trace: src/VX_gather_unit.sv:3:15
											localparam NUM_LANES = _param_8E516_NUM_LANES;
											// Trace: src/VX_gather_unit.sv:4:15
											localparam OUT_BUF = _param_8E516_OUT_BUF;
											// Trace: src/VX_gather_unit.sv:6:5
											wire clk;
											// Trace: src/VX_gather_unit.sv:7:5
											wire reset;
											// Trace: src/VX_gather_unit.sv:8:5
											localparam _mbase_commit_in_if = 0;
											// Trace: src/VX_gather_unit.sv:9:5
											localparam _mbase_commit_out_if = 0;
											// Trace: src/VX_gather_unit.sv:11:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_gather_unit.sv:12:5
											localparam PID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:13:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:14:5
											localparam DATAW = 176;
											// Trace: src/VX_gather_unit.sv:15:5
											localparam DATA_WIS_OFF = 173;
											// Trace: src/VX_gather_unit.sv:16:5
											wire [0:0] commit_in_valid;
											// Trace: src/VX_gather_unit.sv:17:5
											wire [175:0] commit_in_data;
											// Trace: src/VX_gather_unit.sv:18:5
											wire [0:0] commit_in_ready;
											// Trace: src/VX_gather_unit.sv:19:5
											localparam VX_gpu_pkg_ISSUE_ISW = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											wire [0:0] commit_in_isw;
											// Trace: src/VX_gather_unit.sv:20:5
											genvar _gv_i_208;
											for (_gv_i_208 = 0; _gv_i_208 < BLOCK_SIZE; _gv_i_208 = _gv_i_208 + 1) begin : g_commit_in
												localparam i = _gv_i_208;
												// Trace: src/VX_gather_unit.sv:21:9
												assign commit_in_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_commit_if[i + _mbase_commit_in_if].valid;
												// Trace: src/VX_gather_unit.sv:22:9
												assign commit_in_data[i * 176+:176] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_commit_if[i + _mbase_commit_in_if].data;
												// Trace: src/VX_gather_unit.sv:23:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_commit_if[i + _mbase_commit_in_if].ready = commit_in_ready[i];
												if (1) begin : g_commit_in_isw_full
													// Trace: src/VX_gather_unit.sv:31:13
													assign commit_in_isw[i+:1] = sv2v_cast_1_signed(i);
												end
											end
											// Trace: src/VX_gather_unit.sv:34:5
											reg [0:0] commit_out_valid;
											// Trace: src/VX_gather_unit.sv:35:5
											reg [175:0] commit_out_data;
											// Trace: src/VX_gather_unit.sv:36:5
											wire [0:0] commit_out_ready;
											// Trace: src/VX_gather_unit.sv:37:5
											always @(*) begin
												// Trace: src/VX_gather_unit.sv:38:9
												commit_out_valid = 1'sb0;
												// Trace: src/VX_gather_unit.sv:39:9
												begin : sv2v_autoblock_10
													// Trace: src/VX_gather_unit.sv:39:14
													integer i;
													// Trace: src/VX_gather_unit.sv:39:14
													for (i = 0; i < 1; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:40:13
															commit_out_data[i * 176+:176] = 1'sbx;
														end
												end
												begin : sv2v_autoblock_11
													// Trace: src/VX_gather_unit.sv:42:14
													integer i;
													// Trace: src/VX_gather_unit.sv:42:14
													for (i = 0; i < BLOCK_SIZE; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:43:13
															commit_out_valid[commit_in_isw[i+:1]] = commit_in_valid[i];
															// Trace: src/VX_gather_unit.sv:44:13
															commit_out_data[commit_in_isw[i+:1] * 176+:176] = commit_in_data[i * 176+:176];
														end
												end
											end
											// Trace: src/VX_gather_unit.sv:47:5
											genvar _gv_i_209;
											for (_gv_i_209 = 0; _gv_i_209 < BLOCK_SIZE; _gv_i_209 = _gv_i_209 + 1) begin : g_commit_in_ready
												localparam i = _gv_i_209;
												// Trace: src/VX_gather_unit.sv:48:9
												assign commit_in_ready[i] = commit_out_ready[commit_in_isw[i+:1]];
											end
											// Trace: src/VX_gather_unit.sv:50:5
											genvar _gv_i_210;
											for (_gv_i_210 = 0; _gv_i_210 < 1; _gv_i_210 = _gv_i_210 + 1) begin : g_out_bufs
												localparam i = _gv_i_210;
												// Trace: src/VX_gather_unit.sv:51:9
												// expanded interface instance: commit_tmp_if
												localparam _param_C9958_NUM_LANES = NUM_LANES;
												if (1) begin : commit_tmp_if
													// Trace: src/VX_commit_if.sv:2:15
													localparam NUM_LANES = _param_C9958_NUM_LANES;
													// Trace: src/VX_commit_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_commit_if.sv:5:5
													// removed localparam type data_t
													// Trace: src/VX_commit_if.sv:17:5
													wire valid;
													// Trace: src/VX_commit_if.sv:18:5
													wire [175:0] data;
													// Trace: src/VX_commit_if.sv:19:5
													wire ready;
													// Trace: src/VX_commit_if.sv:20:5
													// Trace: src/VX_commit_if.sv:25:5
												end
												// Trace: src/VX_gather_unit.sv:54:9
												VX_elastic_buffer #(
													.DATAW(DATAW),
													.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
													.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
												) out_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(commit_out_valid[i]),
													.ready_in(commit_out_ready[i]),
													.data_in(commit_out_data[i * 176+:176]),
													.data_out(commit_tmp_if.data),
													.valid_out(commit_tmp_if.valid),
													.ready_out(commit_tmp_if.ready)
												);
												// Trace: src/VX_gather_unit.sv:68:9
												wire [3:0] commit_tmask_w;
												// Trace: src/VX_gather_unit.sv:69:9
												wire [127:0] commit_data_w;
												if (1) begin : g_commit_data_no_pid
													// Trace: src/VX_gather_unit.sv:80:13
													assign commit_tmask_w = commit_tmp_if.data[172-:4];
													// Trace: src/VX_gather_unit.sv:81:13
													assign commit_data_w = commit_tmp_if.data[130-:128];
												end
												// Trace: src/VX_gather_unit.sv:83:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].valid = commit_tmp_if.valid;
												// Trace: src/VX_gather_unit.sv:84:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].data = {commit_tmp_if.data[175], commit_tmp_if.data[174-:2], commit_tmask_w, commit_tmp_if.data[168-:31], commit_tmp_if.data[137], commit_tmp_if.data[136-:6], commit_data_w, 1'b0, commit_tmp_if.data[1], commit_tmp_if.data[0]};
												// Trace: src/VX_gather_unit.sv:96:9
												assign commit_tmp_if.ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].ready;
											end
										end
										assign gather_unit.clk = clk;
										assign gather_unit.reset = reset;
									end
									assign alu_unit.clk = clk;
									assign alu_unit.reset = reset;
									// Trace: src/VX_execute.sv:27:5
									// expanded module instance: lsu_unit
									localparam _bbase_54826_dispatch_if = 1;
									localparam _bbase_54826_commit_if = 1;
									localparam _bbase_54826_lsu_mem_if = 0;
									localparam _param_54826_INSTANCE_ID = "";
									if (1) begin : lsu_unit
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_lsu_unit.sv:2:16
										localparam INSTANCE_ID = _param_54826_INSTANCE_ID;
										// Trace: src/VX_lsu_unit.sv:4:5
										wire clk;
										// Trace: src/VX_lsu_unit.sv:5:5
										wire reset;
										// Trace: src/VX_lsu_unit.sv:6:5
										localparam _mbase_dispatch_if = 1;
										// Trace: src/VX_lsu_unit.sv:7:5
										localparam _mbase_commit_if = 1;
										// Trace: src/VX_lsu_unit.sv:8:5
										localparam _mbase_lsu_mem_if = 0;
										// Trace: src/VX_lsu_unit.sv:10:5
										localparam BLOCK_SIZE = 1;
										// Trace: src/VX_lsu_unit.sv:11:5
										localparam NUM_LANES = 4;
										// Trace: src/VX_lsu_unit.sv:13:5
										// expanded interface instance: per_block_execute_if
										localparam _param_E2592_NUM_LANES = NUM_LANES;
										genvar _arr_E2592;
										for (_arr_E2592 = 0; _arr_E2592 <= 0; _arr_E2592 = _arr_E2592 + 1) begin : per_block_execute_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_execute_if.sv:2:15
											localparam NUM_LANES = _param_E2592_NUM_LANES;
											// Trace: src/VX_execute_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_execute_if.sv:5:5
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_execute_if.sv:22:5
											wire valid;
											// Trace: src/VX_execute_if.sv:23:5
											wire [474:0] data;
											// Trace: src/VX_execute_if.sv:24:5
											wire ready;
											// Trace: src/VX_execute_if.sv:25:5
											// Trace: src/VX_execute_if.sv:30:5
										end
										// Trace: src/VX_lsu_unit.sv:16:5
										// expanded module instance: dispatch_unit
										localparam _bbase_2E16E_dispatch_if = 1;
										localparam _bbase_2E16E_execute_if = 0;
										localparam _param_2E16E_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_2E16E_NUM_LANES = NUM_LANES;
										localparam _param_2E16E_OUT_BUF = 3;
										if (1) begin : dispatch_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_dispatch_unit.sv:2:15
											localparam BLOCK_SIZE = _param_2E16E_BLOCK_SIZE;
											// Trace: src/VX_dispatch_unit.sv:3:15
											localparam NUM_LANES = _param_2E16E_NUM_LANES;
											// Trace: src/VX_dispatch_unit.sv:4:15
											localparam OUT_BUF = _param_2E16E_OUT_BUF;
											// Trace: src/VX_dispatch_unit.sv:5:15
											localparam MAX_FANOUT = 8;
											// Trace: src/VX_dispatch_unit.sv:7:5
											wire clk;
											// Trace: src/VX_dispatch_unit.sv:8:5
											wire reset;
											// Trace: src/VX_dispatch_unit.sv:9:5
											localparam _mbase_dispatch_if = 1;
											// Trace: src/VX_dispatch_unit.sv:10:5
											localparam _mbase_execute_if = 0;
											// Trace: src/VX_dispatch_unit.sv:12:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:13:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_dispatch_unit.sv:14:5
											localparam PID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:15:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:16:5
											localparam BATCH_COUNT = 1;
											// Trace: src/VX_dispatch_unit.sv:17:5
											localparam BATCH_COUNT_W = 1;
											// Trace: src/VX_dispatch_unit.sv:18:5
											localparam ISSUE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:19:5
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											localparam VX_gpu_pkg_ISSUE_WIS = 2;
											localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											localparam IN_DATAW = 472;
											// Trace: src/VX_dispatch_unit.sv:20:5
											localparam OUT_DATAW = 475;
											// Trace: src/VX_dispatch_unit.sv:21:5
											localparam FANOUT_ENABLE = 1'd0;
											// Trace: src/VX_dispatch_unit.sv:22:5
											localparam DATA_TMASK_OFF = 465;
											// Trace: src/VX_dispatch_unit.sv:23:5
											localparam DATA_REGS_OFF = 0;
											// Trace: src/VX_dispatch_unit.sv:24:5
											wire [0:0] dispatch_valid;
											// Trace: src/VX_dispatch_unit.sv:25:5
											wire [471:0] dispatch_data;
											// Trace: src/VX_dispatch_unit.sv:26:5
											wire [0:0] dispatch_ready;
											// Trace: src/VX_dispatch_unit.sv:27:5
											genvar _gv_i_96;
											for (_gv_i_96 = 0; _gv_i_96 < 1; _gv_i_96 = _gv_i_96 + 1) begin : g_dispatch_data
												localparam i = _gv_i_96;
												// Trace: src/VX_dispatch_unit.sv:28:9
												assign dispatch_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].valid;
												// Trace: src/VX_dispatch_unit.sv:29:9
												assign dispatch_data[i * 472+:472] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].data;
												// Trace: src/VX_dispatch_unit.sv:30:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].ready = dispatch_ready[i];
											end
											// Trace: src/VX_dispatch_unit.sv:32:5
											wire [0:0] block_ready;
											// Trace: src/VX_dispatch_unit.sv:33:5
											wire [3:0] block_tmask;
											// Trace: src/VX_dispatch_unit.sv:34:5
											wire [383:0] block_regs;
											// Trace: src/VX_dispatch_unit.sv:35:5
											wire [0:0] block_pid;
											// Trace: src/VX_dispatch_unit.sv:36:5
											wire [0:0] block_sop;
											// Trace: src/VX_dispatch_unit.sv:37:5
											wire [0:0] block_eop;
											// Trace: src/VX_dispatch_unit.sv:38:5
											wire [0:0] block_done;
											// Trace: src/VX_dispatch_unit.sv:39:5
											wire batch_done = &block_done;
											// Trace: src/VX_dispatch_unit.sv:40:5
											wire [0:0] batch_idx;
											// Trace: src/VX_dispatch_unit.sv:41:5
											if (1) begin : g_batch_idx_0
												// Trace: src/VX_dispatch_unit.sv:67:9
												assign batch_idx = 0;
											end
											// Trace: src/VX_dispatch_unit.sv:69:5
											wire [0:0] issue_indices;
											// Trace: src/VX_dispatch_unit.sv:70:5
											genvar _gv_block_idx_2;
											for (_gv_block_idx_2 = 0; _gv_block_idx_2 < BLOCK_SIZE; _gv_block_idx_2 = _gv_block_idx_2 + 1) begin : g_issue_indices
												localparam block_idx = _gv_block_idx_2;
												// Trace: src/VX_dispatch_unit.sv:71:9
												assign issue_indices[block_idx+:1] = sv2v_cast_1(batch_idx * BLOCK_SIZE) + sv2v_cast_1_signed(block_idx);
											end
											// Trace: src/VX_dispatch_unit.sv:73:5
											genvar _gv_block_idx_3;
											localparam VX_gpu_pkg_ISSUE_ISW = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											function [1:0] VX_gpu_pkg_wis_to_wid;
												// Trace: src/VX_gpu_pkg.sv:151:9
												input reg [1:0] wis;
												// Trace: src/VX_gpu_pkg.sv:152:9
												input reg [0:0] isw;
												// Trace: src/VX_gpu_pkg.sv:154:9
												begin
													// Trace: src/VX_gpu_pkg.sv:157:13
													VX_gpu_pkg_wis_to_wid = wis;
												end
											endfunction
											for (_gv_block_idx_3 = 0; _gv_block_idx_3 < BLOCK_SIZE; _gv_block_idx_3 = _gv_block_idx_3 + 1) begin : g_blocks
												localparam block_idx = _gv_block_idx_3;
												// Trace: src/VX_dispatch_unit.sv:74:9
												wire [0:0] issue_idx = issue_indices[block_idx+:1];
												// Trace: src/VX_dispatch_unit.sv:75:9
												wire valid_p;
												wire ready_p;
												if (1) begin : g_full_threads
													// Trace: src/VX_dispatch_unit.sv:168:13
													assign valid_p = dispatch_valid[issue_idx];
													// Trace: src/VX_dispatch_unit.sv:169:13
													assign block_tmask[block_idx * 4+:4] = dispatch_data[(issue_idx * 472) + DATA_TMASK_OFF+:4];
													// Trace: src/VX_dispatch_unit.sv:170:13
													assign block_regs[32 * ((block_idx * 3) * 4)+:128] = dispatch_data[(issue_idx * 472) + 256+:128];
													// Trace: src/VX_dispatch_unit.sv:171:13
													assign block_regs[32 * (((block_idx * 3) + 1) * 4)+:128] = dispatch_data[(issue_idx * 472) + 128+:128];
													// Trace: src/VX_dispatch_unit.sv:172:13
													assign block_regs[32 * (((block_idx * 3) + 2) * 4)+:128] = dispatch_data[issue_idx * 472+:128];
													// Trace: src/VX_dispatch_unit.sv:173:13
													assign block_pid[block_idx+:1] = 1'sb0;
													// Trace: src/VX_dispatch_unit.sv:174:13
													assign block_sop[block_idx] = 1'b1;
													// Trace: src/VX_dispatch_unit.sv:175:13
													assign block_eop[block_idx] = 1'b1;
													// Trace: src/VX_dispatch_unit.sv:176:13
													assign block_ready[block_idx] = ready_p;
													// Trace: src/VX_dispatch_unit.sv:177:13
													assign block_done[block_idx] = ready_p || ~valid_p;
												end
												// Trace: src/VX_dispatch_unit.sv:179:9
												wire [0:0] isw;
												if (1) begin : g_isw
													// Trace: src/VX_dispatch_unit.sv:187:13
													assign isw = block_idx;
												end
												// Trace: src/VX_dispatch_unit.sv:189:9
												wire [1:0] block_wid = VX_gpu_pkg_wis_to_wid(dispatch_data[(issue_idx * 472) + 469+:VX_gpu_pkg_ISSUE_WIS_W], isw);
												// Trace: src/VX_dispatch_unit.sv:190:9
												wire [474:0] execute_data;
												reg [474:0] execute_data_w;
												// Trace: src/VX_dispatch_unit.sv:191:9
												VX_elastic_buffer #(
													.DATAW(OUT_DATAW),
													.SIZE(2),
													.OUT_REG(1)
												) buf_out(
													.clk(clk),
													.reset(reset),
													.valid_in(valid_p),
													.ready_in(ready_p),
													.data_in({dispatch_data[(issue_idx * 472) + 471-:1], block_wid, block_tmask[block_idx * 4+:4], dispatch_data[(issue_idx * 472) + 464-:81], block_regs[32 * ((block_idx * 3) * 4)+:128], block_regs[32 * (((block_idx * 3) + 1) * 4)+:128], block_regs[32 * (((block_idx * 3) + 2) * 4)+:128], block_pid[block_idx+:1], block_sop[block_idx], block_eop[block_idx]}),
													.data_out(execute_data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[block_idx + _mbase_execute_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[block_idx + _mbase_execute_if].ready)
												);
												if (1) begin : g_execute_data_w_full
													// Trace: src/VX_dispatch_unit.sv:218:13
													always @(*) begin
														// Trace: src/VX_dispatch_unit.sv:219:17
														execute_data_w = execute_data;
														// Trace: src/VX_dispatch_unit.sv:220:17
														execute_data_w[2:0] = 3'b011;
													end
												end
												// Trace: src/VX_dispatch_unit.sv:223:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[block_idx + _mbase_execute_if].data = execute_data_w;
											end
											// Trace: src/VX_dispatch_unit.sv:225:5
											reg [0:0] ready_in;
											// Trace: src/VX_dispatch_unit.sv:226:5
											always @(*) begin
												// Trace: src/VX_dispatch_unit.sv:227:9
												ready_in = 0;
												// Trace: src/VX_dispatch_unit.sv:228:9
												begin : sv2v_autoblock_12
													// Trace: src/VX_dispatch_unit.sv:228:14
													integer block_idx;
													// Trace: src/VX_dispatch_unit.sv:228:14
													for (block_idx = 0; block_idx < BLOCK_SIZE; block_idx = block_idx + 1)
														begin
															// Trace: src/VX_dispatch_unit.sv:229:13
															ready_in[issue_indices[block_idx+:1]] = block_ready[block_idx] && block_eop[block_idx];
														end
												end
											end
											// Trace: src/VX_dispatch_unit.sv:232:5
											assign dispatch_ready = ready_in;
										end
										assign dispatch_unit.clk = clk;
										assign dispatch_unit.reset = reset;
										// Trace: src/VX_lsu_unit.sv:26:5
										// expanded interface instance: per_block_commit_if
										localparam _param_98792_NUM_LANES = NUM_LANES;
										genvar _arr_98792;
										for (_arr_98792 = 0; _arr_98792 <= 0; _arr_98792 = _arr_98792 + 1) begin : per_block_commit_if
											// Trace: src/VX_commit_if.sv:2:15
											localparam NUM_LANES = _param_98792_NUM_LANES;
											// Trace: src/VX_commit_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_commit_if.sv:5:5
											// removed localparam type data_t
											// Trace: src/VX_commit_if.sv:17:5
											wire valid;
											// Trace: src/VX_commit_if.sv:18:5
											wire [175:0] data;
											// Trace: src/VX_commit_if.sv:19:5
											wire ready;
											// Trace: src/VX_commit_if.sv:20:5
											// Trace: src/VX_commit_if.sv:25:5
										end
										// Trace: src/VX_lsu_unit.sv:29:5
										genvar _gv_block_idx_1;
										for (_gv_block_idx_1 = 0; _gv_block_idx_1 < BLOCK_SIZE; _gv_block_idx_1 = _gv_block_idx_1 + 1) begin : g_slices
											localparam block_idx = _gv_block_idx_1;
											// Trace: src/VX_lsu_unit.sv:30:9
											// expanded module instance: lsu_slice
											localparam _bbase_DE6D2_execute_if = block_idx;
											localparam _bbase_DE6D2_commit_if = block_idx;
											localparam _bbase_DE6D2_lsu_mem_if = block_idx + _mbase_lsu_mem_if;
											localparam _param_DE6D2_INSTANCE_ID = "";
											if (1) begin : lsu_slice
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_lsu_slice.sv:2:16
												localparam INSTANCE_ID = _param_DE6D2_INSTANCE_ID;
												// Trace: src/VX_lsu_slice.sv:4:5
												wire clk;
												// Trace: src/VX_lsu_slice.sv:5:5
												wire reset;
												// Trace: src/VX_lsu_slice.sv:6:5
												localparam _mbase_execute_if = _bbase_DE6D2_execute_if;
												// Trace: src/VX_lsu_slice.sv:7:5
												localparam _mbase_commit_if = _bbase_DE6D2_commit_if;
												// Trace: src/VX_lsu_slice.sv:8:5
												localparam _mbase_lsu_mem_if = _bbase_DE6D2_lsu_mem_if;
												// Trace: src/VX_lsu_slice.sv:10:5
												localparam NUM_LANES = 4;
												// Trace: src/VX_lsu_slice.sv:11:5
												localparam PID_BITS = 0;
												// Trace: src/VX_lsu_slice.sv:12:5
												localparam PID_WIDTH = 1;
												// Trace: src/VX_lsu_slice.sv:13:5
												localparam RSP_ARB_DATAW = 176;
												// Trace: src/VX_lsu_slice.sv:14:5
												localparam LSUQ_SIZEW = 1;
												// Trace: src/VX_lsu_slice.sv:15:5
												localparam VX_gpu_pkg_LSU_WORD_SIZE = 4;
												localparam REQ_ASHIFT = 2;
												// Trace: src/VX_lsu_slice.sv:16:5
												localparam MEM_ASHIFT = 6;
												// Trace: src/VX_lsu_slice.sv:17:5
												localparam MEM_ADDRW = 26;
												// Trace: src/VX_lsu_slice.sv:18:5
												localparam TAG_ID_WIDTH = 55;
												// Trace: src/VX_lsu_slice.sv:19:5
												localparam TAG_WIDTH = 56;
												// Trace: src/VX_lsu_slice.sv:20:5
												// expanded interface instance: commit_rsp_if
												localparam _param_1FB24_NUM_LANES = NUM_LANES;
												if (1) begin : commit_rsp_if
													// Trace: src/VX_commit_if.sv:2:15
													localparam NUM_LANES = _param_1FB24_NUM_LANES;
													// Trace: src/VX_commit_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_commit_if.sv:5:5
													// removed localparam type data_t
													// Trace: src/VX_commit_if.sv:17:5
													wire valid;
													// Trace: src/VX_commit_if.sv:18:5
													wire [175:0] data;
													// Trace: src/VX_commit_if.sv:19:5
													wire ready;
													// Trace: src/VX_commit_if.sv:20:5
													// Trace: src/VX_commit_if.sv:25:5
												end
												// Trace: src/VX_lsu_slice.sv:23:5
												// expanded interface instance: commit_no_rsp_if
												localparam _param_23ED7_NUM_LANES = NUM_LANES;
												if (1) begin : commit_no_rsp_if
													// Trace: src/VX_commit_if.sv:2:15
													localparam NUM_LANES = _param_23ED7_NUM_LANES;
													// Trace: src/VX_commit_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_commit_if.sv:5:5
													// removed localparam type data_t
													// Trace: src/VX_commit_if.sv:17:5
													wire valid;
													// Trace: src/VX_commit_if.sv:18:5
													wire [175:0] data;
													// Trace: src/VX_commit_if.sv:19:5
													wire ready;
													// Trace: src/VX_commit_if.sv:20:5
													// Trace: src/VX_commit_if.sv:25:5
												end
												// Trace: src/VX_lsu_slice.sv:26:5
												wire req_is_fence;
												wire rsp_is_fence;
												// Trace: src/VX_lsu_slice.sv:27:5
												wire [127:0] full_addr;
												// Trace: src/VX_lsu_slice.sv:28:5
												genvar _gv_i_51;
												for (_gv_i_51 = 0; _gv_i_51 < NUM_LANES; _gv_i_51 = _gv_i_51 + 1) begin : g_full_addr
													localparam i = _gv_i_51;
													// Trace: src/VX_lsu_slice.sv:29:9
													assign full_addr[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[259 + (i * 32)+:32] + {{21 {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[407]}}, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[406:396]};
												end
												// Trace: src/VX_lsu_slice.sv:31:5
												wire [11:0] mem_req_flags;
												// Trace: src/VX_lsu_slice.sv:32:5
												genvar _gv_i_52;
												for (_gv_i_52 = 0; _gv_i_52 < NUM_LANES; _gv_i_52 = _gv_i_52 + 1) begin : g_mem_req_flags
													localparam i = _gv_i_52;
													// Trace: src/VX_lsu_slice.sv:33:9
													wire [25:0] block_addr = full_addr[(i * 32) + MEM_ASHIFT+:MEM_ADDRW];
													// Trace: src/VX_lsu_slice.sv:34:9
													wire [25:0] io_addr_start = sv2v_cast_26(32'h00000040 >> MEM_ASHIFT);
													// Trace: src/VX_lsu_slice.sv:35:9
													wire [25:0] io_addr_end = sv2v_cast_26(32'h00010000 >> MEM_ASHIFT);
													// Trace: src/VX_lsu_slice.sv:36:9
													assign mem_req_flags[i * 3] = req_is_fence;
													// Trace: src/VX_lsu_slice.sv:37:9
													assign mem_req_flags[(i * 3) + 1] = (block_addr >= io_addr_start) && (block_addr < io_addr_end);
													// Trace: src/VX_lsu_slice.sv:38:9
													wire [25:0] lmem_addr_start = sv2v_cast_26(32'hffff0000 >> MEM_ASHIFT);
													// Trace: src/VX_lsu_slice.sv:39:9
													wire [25:0] lmem_addr_end = sv2v_cast_26((32'hffff0000 + 32'sd16384) >> MEM_ASHIFT);
													// Trace: src/VX_lsu_slice.sv:40:9
													assign mem_req_flags[(i * 3) + 2] = (block_addr >= lmem_addr_start) && (block_addr < lmem_addr_end);
												end
												// Trace: src/VX_lsu_slice.sv:42:5
												wire mem_req_valid;
												// Trace: src/VX_lsu_slice.sv:43:5
												wire [3:0] mem_req_mask;
												// Trace: src/VX_lsu_slice.sv:44:5
												wire mem_req_rw;
												// Trace: src/VX_lsu_slice.sv:45:5
												localparam VX_gpu_pkg_LSU_ADDR_WIDTH = 30;
												wire [119:0] mem_req_addr;
												// Trace: src/VX_lsu_slice.sv:46:5
												wire [15:0] mem_req_byteen;
												// Trace: src/VX_lsu_slice.sv:47:5
												reg [127:0] mem_req_data;
												// Trace: src/VX_lsu_slice.sv:48:5
												wire [55:0] mem_req_tag;
												// Trace: src/VX_lsu_slice.sv:49:5
												wire mem_req_ready;
												// Trace: src/VX_lsu_slice.sv:50:5
												wire mem_rsp_valid;
												// Trace: src/VX_lsu_slice.sv:51:5
												wire [3:0] mem_rsp_mask;
												// Trace: src/VX_lsu_slice.sv:52:5
												wire [127:0] mem_rsp_data;
												// Trace: src/VX_lsu_slice.sv:53:5
												wire [55:0] mem_rsp_tag;
												// Trace: src/VX_lsu_slice.sv:54:5
												wire mem_rsp_sop;
												// Trace: src/VX_lsu_slice.sv:55:5
												wire mem_rsp_eop;
												// Trace: src/VX_lsu_slice.sv:56:5
												wire mem_rsp_ready;
												// Trace: src/VX_lsu_slice.sv:57:5
												wire mem_req_fire = mem_req_valid && mem_req_ready;
												// Trace: src/VX_lsu_slice.sv:58:5
												wire mem_rsp_fire = mem_rsp_valid && mem_rsp_ready;
												// Trace: src/VX_lsu_slice.sv:59:5
												wire mem_rsp_sop_pkt;
												wire mem_rsp_eop_pkt;
												// Trace: src/VX_lsu_slice.sv:60:5
												wire no_rsp_buf_valid;
												wire no_rsp_buf_ready;
												// Trace: src/VX_lsu_slice.sv:61:5
												reg fence_lock;
												// Trace: src/VX_lsu_slice.sv:62:5
												assign req_is_fence = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[436:435] == 3;
												// Trace: src/VX_lsu_slice.sv:63:5
												always @(posedge clk)
													// Trace: src/VX_lsu_slice.sv:64:9
													if (reset)
														// Trace: src/VX_lsu_slice.sv:65:13
														fence_lock <= 0;
													else begin
														// Trace: src/VX_lsu_slice.sv:67:13
														if ((mem_req_fire && req_is_fence) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[0])
															// Trace: src/VX_lsu_slice.sv:68:17
															fence_lock <= 1;
														if ((mem_rsp_fire && rsp_is_fence) && mem_rsp_eop_pkt)
															// Trace: src/VX_lsu_slice.sv:71:17
															fence_lock <= 0;
													end
												// Trace: src/VX_lsu_slice.sv:75:5
												wire req_skip = req_is_fence && ~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[0];
												// Trace: src/VX_lsu_slice.sv:76:5
												wire no_rsp_buf_enable = (mem_req_rw && ~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[395]) || req_skip;
												// Trace: src/VX_lsu_slice.sv:77:5
												assign mem_req_valid = ((Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].valid && ~req_skip) && ~(no_rsp_buf_enable && ~no_rsp_buf_ready)) && ~fence_lock;
												// Trace: src/VX_lsu_slice.sv:81:5
												assign no_rsp_buf_valid = ((Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].valid && no_rsp_buf_enable) && (req_skip || mem_req_ready)) && ~fence_lock;
												// Trace: src/VX_lsu_slice.sv:85:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].ready = ((mem_req_ready || req_skip) && ~(no_rsp_buf_enable && ~no_rsp_buf_ready)) && ~fence_lock;
												// Trace: src/VX_lsu_slice.sv:88:5
												assign mem_req_mask = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[471-:4];
												// Trace: src/VX_lsu_slice.sv:89:5
												assign mem_req_rw = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[409];
												// Trace: src/VX_lsu_slice.sv:90:5
												wire [7:0] req_align;
												// Trace: src/VX_lsu_slice.sv:91:5
												genvar _gv_i_53;
												for (_gv_i_53 = 0; _gv_i_53 < NUM_LANES; _gv_i_53 = _gv_i_53 + 1) begin : g_mem_req_addr
													localparam i = _gv_i_53;
													// Trace: src/VX_lsu_slice.sv:92:9
													assign req_align[i * 2+:2] = full_addr[(i * 32) + 1-:2];
													// Trace: src/VX_lsu_slice.sv:93:9
													assign mem_req_addr[i * 30+:30] = full_addr[(i * 32) + 31-:30];
												end
												// Trace: src/VX_lsu_slice.sv:95:5
												genvar _gv_i_54;
												for (_gv_i_54 = 0; _gv_i_54 < NUM_LANES; _gv_i_54 = _gv_i_54 + 1) begin : g_mem_req_byteen_w
													localparam i = _gv_i_54;
													// Trace: src/VX_lsu_slice.sv:96:9
													reg [3:0] mem_req_byteen_w;
													// Trace: src/VX_lsu_slice.sv:97:9
													always @(*) begin
														// Trace: src/VX_lsu_slice.sv:98:13
														mem_req_byteen_w = 1'sb0;
														// Trace: src/VX_lsu_slice.sv:99:13
														case (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[434:433])
															0:
																// Trace: src/VX_lsu_slice.sv:101:21
																mem_req_byteen_w[req_align[i * 2+:2]] = 1'b1;
															1: begin
																// Trace: src/VX_lsu_slice.sv:104:21
																mem_req_byteen_w[{req_align[(i * 2) + 1-:1], 1'b0}] = 1'b1;
																// Trace: src/VX_lsu_slice.sv:105:21
																mem_req_byteen_w[{req_align[(i * 2) + 1-:1], 1'b1}] = 1'b1;
															end
															default:
																// Trace: src/VX_lsu_slice.sv:107:27
																mem_req_byteen_w = {VX_gpu_pkg_LSU_WORD_SIZE {1'b1}};
														endcase
													end
													// Trace: src/VX_lsu_slice.sv:110:9
													assign mem_req_byteen[i * 4+:4] = mem_req_byteen_w;
												end
												// Trace: src/VX_lsu_slice.sv:112:5
												genvar _gv_i_55;
												for (_gv_i_55 = 0; _gv_i_55 < NUM_LANES; _gv_i_55 = _gv_i_55 + 1) begin : g_missalign
													localparam i = _gv_i_55;
													// Trace: src/VX_lsu_slice.sv:113:9
													wire lsu_req_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].ready;
												end
												// Trace: src/VX_lsu_slice.sv:115:5
												genvar _gv_i_56;
												for (_gv_i_56 = 0; _gv_i_56 < NUM_LANES; _gv_i_56 = _gv_i_56 + 1) begin : g_mem_req_data
													localparam i = _gv_i_56;
													// Trace: src/VX_lsu_slice.sv:116:9
													always @(*) begin
														// Trace: src/VX_lsu_slice.sv:117:13
														mem_req_data[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[131 + (i * 32)+:32];
														// Trace: src/VX_lsu_slice.sv:118:13
														case (req_align[i * 2+:2])
															1:
																// Trace: src/VX_lsu_slice.sv:119:20
																mem_req_data[(i * 32) + 31-:24] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[131 + ((i * 32) + 23)-:24];
															2:
																// Trace: src/VX_lsu_slice.sv:120:20
																mem_req_data[(i * 32) + 31-:16] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[131 + ((i * 32) + 15)-:16];
															3:
																// Trace: src/VX_lsu_slice.sv:121:20
																mem_req_data[(i * 32) + 31-:8] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[131 + ((i * 32) + 7)-:8];
															default:
																;
														endcase
													end
												end
												// Trace: src/VX_lsu_slice.sv:126:5
												wire [0:0] pkt_waddr;
												wire [0:0] pkt_raddr;
												// Trace: src/VX_lsu_slice.sv:127:5
												if (1) begin : g_no_pids
													// Trace: src/VX_lsu_slice.sv:179:9
													assign pkt_waddr = 0;
													// Trace: src/VX_lsu_slice.sv:180:9
													assign mem_rsp_sop_pkt = mem_rsp_sop;
													// Trace: src/VX_lsu_slice.sv:181:9
													assign mem_rsp_eop_pkt = mem_rsp_eop;
												end
												// Trace: src/VX_lsu_slice.sv:183:5
												assign mem_req_tag = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[474], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[473-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[467-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[395], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[394-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[436-:4], req_align, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[2], pkt_waddr, req_is_fence};
												// Trace: src/VX_lsu_slice.sv:195:5
												wire lsu_mem_req_valid;
												// Trace: src/VX_lsu_slice.sv:196:5
												wire lsu_mem_req_rw;
												// Trace: src/VX_lsu_slice.sv:197:5
												wire [3:0] lsu_mem_req_mask;
												// Trace: src/VX_lsu_slice.sv:198:5
												wire [15:0] lsu_mem_req_byteen;
												// Trace: src/VX_lsu_slice.sv:199:5
												wire [119:0] lsu_mem_req_addr;
												// Trace: src/VX_lsu_slice.sv:200:5
												wire [11:0] lsu_mem_req_flags;
												// Trace: src/VX_lsu_slice.sv:201:5
												wire [127:0] lsu_mem_req_data;
												// Trace: src/VX_lsu_slice.sv:202:5
												localparam VX_gpu_pkg_LSU_MEM_BATCHES = 1;
												localparam VX_gpu_pkg_LSU_TAG_ID_BITS = 1;
												localparam VX_gpu_pkg_LSU_TAG_WIDTH = 2;
												wire [1:0] lsu_mem_req_tag;
												// Trace: src/VX_lsu_slice.sv:203:5
												wire lsu_mem_req_ready;
												// Trace: src/VX_lsu_slice.sv:204:5
												wire lsu_mem_rsp_valid;
												// Trace: src/VX_lsu_slice.sv:205:5
												wire [3:0] lsu_mem_rsp_mask;
												// Trace: src/VX_lsu_slice.sv:206:5
												wire [127:0] lsu_mem_rsp_data;
												// Trace: src/VX_lsu_slice.sv:207:5
												wire [1:0] lsu_mem_rsp_tag;
												// Trace: src/VX_lsu_slice.sv:208:5
												wire lsu_mem_rsp_ready;
												// Trace: src/VX_lsu_slice.sv:209:5
												VX_mem_scheduler #(
													.INSTANCE_ID(""),
													.CORE_REQS(NUM_LANES),
													.MEM_CHANNELS(NUM_LANES),
													.WORD_SIZE(VX_gpu_pkg_LSU_WORD_SIZE),
													.LINE_SIZE(VX_gpu_pkg_LSU_WORD_SIZE),
													.ADDR_WIDTH(VX_gpu_pkg_LSU_ADDR_WIDTH),
													.FLAGS_WIDTH(3),
													.TAG_WIDTH(TAG_WIDTH),
													.CORE_QUEUE_SIZE(2),
													.MEM_QUEUE_SIZE(4),
													.UUID_WIDTH(1),
													.RSP_PARTIAL(1),
													.MEM_OUT_BUF(0),
													.CORE_OUT_BUF(0)
												) mem_scheduler(
													.clk(clk),
													.reset(reset),
													.core_req_valid(mem_req_valid),
													.core_req_rw(mem_req_rw),
													.core_req_mask(mem_req_mask),
													.core_req_byteen(mem_req_byteen),
													.core_req_addr(mem_req_addr),
													.core_req_flags(mem_req_flags),
													.core_req_data(mem_req_data),
													.core_req_tag(mem_req_tag),
													.core_req_ready(mem_req_ready),
													.core_req_empty(),
													.core_req_wr_notify(),
													.core_rsp_valid(mem_rsp_valid),
													.core_rsp_mask(mem_rsp_mask),
													.core_rsp_data(mem_rsp_data),
													.core_rsp_tag(mem_rsp_tag),
													.core_rsp_sop(mem_rsp_sop),
													.core_rsp_eop(mem_rsp_eop),
													.core_rsp_ready(mem_rsp_ready),
													.mem_req_valid(lsu_mem_req_valid),
													.mem_req_rw(lsu_mem_req_rw),
													.mem_req_mask(lsu_mem_req_mask),
													.mem_req_byteen(lsu_mem_req_byteen),
													.mem_req_addr(lsu_mem_req_addr),
													.mem_req_flags(lsu_mem_req_flags),
													.mem_req_data(lsu_mem_req_data),
													.mem_req_tag(lsu_mem_req_tag),
													.mem_req_ready(lsu_mem_req_ready),
													.mem_rsp_valid(lsu_mem_rsp_valid),
													.mem_rsp_mask(lsu_mem_rsp_mask),
													.mem_rsp_data(lsu_mem_rsp_data),
													.mem_rsp_tag(lsu_mem_rsp_tag),
													.mem_rsp_ready(lsu_mem_rsp_ready)
												);
												// Trace: src/VX_lsu_slice.sv:260:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_valid = lsu_mem_req_valid;
												// Trace: src/VX_lsu_slice.sv:261:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[282-:4] = lsu_mem_req_mask;
												// Trace: src/VX_lsu_slice.sv:262:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[278] = lsu_mem_req_rw;
												// Trace: src/VX_lsu_slice.sv:263:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[29-:16] = lsu_mem_req_byteen;
												// Trace: src/VX_lsu_slice.sv:264:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[277-:120] = lsu_mem_req_addr;
												// Trace: src/VX_lsu_slice.sv:265:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[13-:12] = lsu_mem_req_flags;
												// Trace: src/VX_lsu_slice.sv:266:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[157-:128] = lsu_mem_req_data;
												// Trace: src/VX_lsu_slice.sv:267:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[1-:2] = lsu_mem_req_tag;
												// Trace: src/VX_lsu_slice.sv:268:5
												assign lsu_mem_req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_ready;
												// Trace: src/VX_lsu_slice.sv:269:5
												assign lsu_mem_rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_valid;
												// Trace: src/VX_lsu_slice.sv:270:5
												assign lsu_mem_rsp_mask = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_data[133-:4];
												// Trace: src/VX_lsu_slice.sv:271:5
												assign lsu_mem_rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_data[129-:128];
												// Trace: src/VX_lsu_slice.sv:272:5
												assign lsu_mem_rsp_tag = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_data[1-:2];
												// Trace: src/VX_lsu_slice.sv:273:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_ready = lsu_mem_rsp_ready;
												// Trace: src/VX_lsu_slice.sv:274:5
												wire [0:0] rsp_uuid;
												// Trace: src/VX_lsu_slice.sv:275:5
												wire [1:0] rsp_wid;
												// Trace: src/VX_lsu_slice.sv:276:5
												wire [30:0] rsp_pc;
												// Trace: src/VX_lsu_slice.sv:277:5
												wire rsp_wb;
												// Trace: src/VX_lsu_slice.sv:278:5
												wire [5:0] rsp_rd;
												// Trace: src/VX_lsu_slice.sv:279:5
												wire [3:0] rsp_op_type;
												// Trace: src/VX_lsu_slice.sv:280:5
												wire [7:0] rsp_align;
												// Trace: src/VX_lsu_slice.sv:281:5
												wire [0:0] rsp_pid;
												// Trace: src/VX_lsu_slice.sv:282:5
												assign {rsp_uuid, rsp_wid, rsp_pc, rsp_wb, rsp_rd, rsp_op_type, rsp_align, rsp_pid, pkt_raddr, rsp_is_fence} = mem_rsp_tag;
												// Trace: src/VX_lsu_slice.sv:294:5
												reg [127:0] rsp_data;
												// Trace: src/VX_lsu_slice.sv:295:5
												genvar _gv_i_57;
												for (_gv_i_57 = 0; _gv_i_57 < NUM_LANES; _gv_i_57 = _gv_i_57 + 1) begin : g_rsp_data
													localparam i = _gv_i_57;
													// Trace: src/VX_lsu_slice.sv:296:9
													wire [31:0] rsp_data32 = mem_rsp_data[i * 32+:32];
													// Trace: src/VX_lsu_slice.sv:297:9
													wire [15:0] rsp_data16 = (rsp_align[(i * 2) + 1] ? rsp_data32[31:16] : rsp_data32[15:0]);
													// Trace: src/VX_lsu_slice.sv:298:9
													wire [7:0] rsp_data8 = (rsp_align[i * 2] ? rsp_data16[15:8] : rsp_data16[7:0]);
													// Trace: src/VX_lsu_slice.sv:299:9
													always @(*)
														// Trace: src/VX_lsu_slice.sv:300:13
														case (rsp_op_type[2:0])
															3'b000:
																// Trace: src/VX_lsu_slice.sv:301:22
																rsp_data[i * 32+:32] = sv2v_cast_32_signed($signed(rsp_data8));
															3'b001:
																// Trace: src/VX_lsu_slice.sv:302:22
																rsp_data[i * 32+:32] = sv2v_cast_32_signed($signed(rsp_data16));
															3'b100:
																// Trace: src/VX_lsu_slice.sv:303:21
																rsp_data[i * 32+:32] = sv2v_cast_32($unsigned(rsp_data8));
															3'b101:
																// Trace: src/VX_lsu_slice.sv:304:21
																rsp_data[i * 32+:32] = sv2v_cast_32($unsigned(rsp_data16));
															3'b010:
																// Trace: src/VX_lsu_slice.sv:305:22
																rsp_data[i * 32+:32] = sv2v_cast_32_signed($signed(rsp_data32));
															default:
																// Trace: src/VX_lsu_slice.sv:306:22
																rsp_data[i * 32+:32] = 1'sbx;
														endcase
												end
												// Trace: src/VX_lsu_slice.sv:310:5
												VX_elastic_buffer #(
													.DATAW(176),
													.SIZE(2)
												) rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_rsp_valid),
													.ready_in(mem_rsp_ready),
													.data_in({rsp_uuid, rsp_wid, mem_rsp_mask, rsp_pc, rsp_wb, rsp_rd, rsp_data, rsp_pid, mem_rsp_sop_pkt, mem_rsp_eop_pkt}),
													.data_out({commit_rsp_if.data[175], commit_rsp_if.data[174-:2], commit_rsp_if.data[172-:4], commit_rsp_if.data[168-:31], commit_rsp_if.data[137], commit_rsp_if.data[136-:6], commit_rsp_if.data[130-:128], commit_rsp_if.data[2], commit_rsp_if.data[1], commit_rsp_if.data[0]}),
													.valid_out(commit_rsp_if.valid),
													.ready_out(commit_rsp_if.ready)
												);
												// Trace: src/VX_lsu_slice.sv:323:5
												VX_elastic_buffer #(
													.DATAW(41),
													.SIZE(2)
												) no_rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(no_rsp_buf_valid),
													.ready_in(no_rsp_buf_ready),
													.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[474], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[473-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[471-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[467-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[0]}),
													.data_out({commit_no_rsp_if.data[175], commit_no_rsp_if.data[174-:2], commit_no_rsp_if.data[172-:4], commit_no_rsp_if.data[168-:31], commit_no_rsp_if.data[2], commit_no_rsp_if.data[1], commit_no_rsp_if.data[0]}),
													.valid_out(commit_no_rsp_if.valid),
													.ready_out(commit_no_rsp_if.ready)
												);
												// Trace: src/VX_lsu_slice.sv:336:5
												assign commit_no_rsp_if.data[136-:6] = 1'sb0;
												// Trace: src/VX_lsu_slice.sv:337:5
												assign commit_no_rsp_if.data[137] = 1'b0;
												// Trace: src/VX_lsu_slice.sv:338:5
												assign commit_no_rsp_if.data[130-:128] = commit_rsp_if.data[130-:128];
												// Trace: src/VX_lsu_slice.sv:339:5
												VX_stream_arb #(
													.NUM_INPUTS(2),
													.DATAW(RSP_ARB_DATAW),
													.ARBITER("P"),
													.OUT_BUF(3)
												) rsp_arb(
													.clk(clk),
													.reset(reset),
													.valid_in({commit_no_rsp_if.valid, commit_rsp_if.valid}),
													.ready_in({commit_no_rsp_if.ready, commit_rsp_if.ready}),
													.data_in({commit_no_rsp_if.data, commit_rsp_if.data}),
													.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_commit_if[_mbase_commit_if].data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_commit_if[_mbase_commit_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_commit_if[_mbase_commit_if].ready),
													.sel_out()
												);
											end
											assign lsu_slice.clk = clk;
											assign lsu_slice.reset = reset;
										end
										// Trace: src/VX_lsu_unit.sv:40:5
										// expanded module instance: gather_unit
										localparam _bbase_8E516_commit_in_if = 0;
										localparam _bbase_8E516_commit_out_if = 1;
										localparam _param_8E516_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_8E516_NUM_LANES = NUM_LANES;
										localparam _param_8E516_OUT_BUF = 3;
										if (1) begin : gather_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_gather_unit.sv:2:15
											localparam BLOCK_SIZE = _param_8E516_BLOCK_SIZE;
											// Trace: src/VX_gather_unit.sv:3:15
											localparam NUM_LANES = _param_8E516_NUM_LANES;
											// Trace: src/VX_gather_unit.sv:4:15
											localparam OUT_BUF = _param_8E516_OUT_BUF;
											// Trace: src/VX_gather_unit.sv:6:5
											wire clk;
											// Trace: src/VX_gather_unit.sv:7:5
											wire reset;
											// Trace: src/VX_gather_unit.sv:8:5
											localparam _mbase_commit_in_if = 0;
											// Trace: src/VX_gather_unit.sv:9:5
											localparam _mbase_commit_out_if = 1;
											// Trace: src/VX_gather_unit.sv:11:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_gather_unit.sv:12:5
											localparam PID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:13:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:14:5
											localparam DATAW = 176;
											// Trace: src/VX_gather_unit.sv:15:5
											localparam DATA_WIS_OFF = 173;
											// Trace: src/VX_gather_unit.sv:16:5
											wire [0:0] commit_in_valid;
											// Trace: src/VX_gather_unit.sv:17:5
											wire [175:0] commit_in_data;
											// Trace: src/VX_gather_unit.sv:18:5
											wire [0:0] commit_in_ready;
											// Trace: src/VX_gather_unit.sv:19:5
											localparam VX_gpu_pkg_ISSUE_ISW = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											wire [0:0] commit_in_isw;
											// Trace: src/VX_gather_unit.sv:20:5
											genvar _gv_i_208;
											for (_gv_i_208 = 0; _gv_i_208 < BLOCK_SIZE; _gv_i_208 = _gv_i_208 + 1) begin : g_commit_in
												localparam i = _gv_i_208;
												// Trace: src/VX_gather_unit.sv:21:9
												assign commit_in_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_commit_if[i + _mbase_commit_in_if].valid;
												// Trace: src/VX_gather_unit.sv:22:9
												assign commit_in_data[i * 176+:176] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_commit_if[i + _mbase_commit_in_if].data;
												// Trace: src/VX_gather_unit.sv:23:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_commit_if[i + _mbase_commit_in_if].ready = commit_in_ready[i];
												if (1) begin : g_commit_in_isw_full
													// Trace: src/VX_gather_unit.sv:31:13
													assign commit_in_isw[i+:1] = sv2v_cast_1_signed(i);
												end
											end
											// Trace: src/VX_gather_unit.sv:34:5
											reg [0:0] commit_out_valid;
											// Trace: src/VX_gather_unit.sv:35:5
											reg [175:0] commit_out_data;
											// Trace: src/VX_gather_unit.sv:36:5
											wire [0:0] commit_out_ready;
											// Trace: src/VX_gather_unit.sv:37:5
											always @(*) begin
												// Trace: src/VX_gather_unit.sv:38:9
												commit_out_valid = 1'sb0;
												// Trace: src/VX_gather_unit.sv:39:9
												begin : sv2v_autoblock_13
													// Trace: src/VX_gather_unit.sv:39:14
													integer i;
													// Trace: src/VX_gather_unit.sv:39:14
													for (i = 0; i < 1; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:40:13
															commit_out_data[i * 176+:176] = 1'sbx;
														end
												end
												begin : sv2v_autoblock_14
													// Trace: src/VX_gather_unit.sv:42:14
													integer i;
													// Trace: src/VX_gather_unit.sv:42:14
													for (i = 0; i < BLOCK_SIZE; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:43:13
															commit_out_valid[commit_in_isw[i+:1]] = commit_in_valid[i];
															// Trace: src/VX_gather_unit.sv:44:13
															commit_out_data[commit_in_isw[i+:1] * 176+:176] = commit_in_data[i * 176+:176];
														end
												end
											end
											// Trace: src/VX_gather_unit.sv:47:5
											genvar _gv_i_209;
											for (_gv_i_209 = 0; _gv_i_209 < BLOCK_SIZE; _gv_i_209 = _gv_i_209 + 1) begin : g_commit_in_ready
												localparam i = _gv_i_209;
												// Trace: src/VX_gather_unit.sv:48:9
												assign commit_in_ready[i] = commit_out_ready[commit_in_isw[i+:1]];
											end
											// Trace: src/VX_gather_unit.sv:50:5
											genvar _gv_i_210;
											for (_gv_i_210 = 0; _gv_i_210 < 1; _gv_i_210 = _gv_i_210 + 1) begin : g_out_bufs
												localparam i = _gv_i_210;
												// Trace: src/VX_gather_unit.sv:51:9
												// expanded interface instance: commit_tmp_if
												localparam _param_C9958_NUM_LANES = NUM_LANES;
												if (1) begin : commit_tmp_if
													// Trace: src/VX_commit_if.sv:2:15
													localparam NUM_LANES = _param_C9958_NUM_LANES;
													// Trace: src/VX_commit_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_commit_if.sv:5:5
													// removed localparam type data_t
													// Trace: src/VX_commit_if.sv:17:5
													wire valid;
													// Trace: src/VX_commit_if.sv:18:5
													wire [175:0] data;
													// Trace: src/VX_commit_if.sv:19:5
													wire ready;
													// Trace: src/VX_commit_if.sv:20:5
													// Trace: src/VX_commit_if.sv:25:5
												end
												// Trace: src/VX_gather_unit.sv:54:9
												VX_elastic_buffer #(
													.DATAW(DATAW),
													.SIZE(2),
													.OUT_REG(1)
												) out_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(commit_out_valid[i]),
													.ready_in(commit_out_ready[i]),
													.data_in(commit_out_data[i * 176+:176]),
													.data_out(commit_tmp_if.data),
													.valid_out(commit_tmp_if.valid),
													.ready_out(commit_tmp_if.ready)
												);
												// Trace: src/VX_gather_unit.sv:68:9
												wire [3:0] commit_tmask_w;
												// Trace: src/VX_gather_unit.sv:69:9
												wire [127:0] commit_data_w;
												if (1) begin : g_commit_data_no_pid
													// Trace: src/VX_gather_unit.sv:80:13
													assign commit_tmask_w = commit_tmp_if.data[172-:4];
													// Trace: src/VX_gather_unit.sv:81:13
													assign commit_data_w = commit_tmp_if.data[130-:128];
												end
												// Trace: src/VX_gather_unit.sv:83:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].valid = commit_tmp_if.valid;
												// Trace: src/VX_gather_unit.sv:84:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].data = {commit_tmp_if.data[175], commit_tmp_if.data[174-:2], commit_tmask_w, commit_tmp_if.data[168-:31], commit_tmp_if.data[137], commit_tmp_if.data[136-:6], commit_data_w, 1'b0, commit_tmp_if.data[1], commit_tmp_if.data[0]};
												// Trace: src/VX_gather_unit.sv:96:9
												assign commit_tmp_if.ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].ready;
											end
										end
										assign gather_unit.clk = clk;
										assign gather_unit.reset = reset;
									end
									assign lsu_unit.clk = clk;
									assign lsu_unit.reset = reset;
									// Trace: src/VX_execute.sv:36:5
									// expanded module instance: fpu_unit
									localparam _bbase_88E44_dispatch_if = 3;
									localparam _bbase_88E44_commit_if = 3;
									localparam _bbase_88E44_fpu_csr_if = 0;
									localparam _param_88E44_INSTANCE_ID = "";
									if (1) begin : fpu_unit
										// removed import VX_fpu_pkg::*;
										// Trace: src/VX_fpu_unit.sv:2:16
										localparam INSTANCE_ID = _param_88E44_INSTANCE_ID;
										// Trace: src/VX_fpu_unit.sv:4:5
										wire clk;
										// Trace: src/VX_fpu_unit.sv:5:5
										wire reset;
										// Trace: src/VX_fpu_unit.sv:6:5
										localparam _mbase_dispatch_if = 3;
										// Trace: src/VX_fpu_unit.sv:7:5
										localparam _mbase_commit_if = 3;
										// Trace: src/VX_fpu_unit.sv:8:5
										localparam _mbase_fpu_csr_if = 0;
										// Trace: src/VX_fpu_unit.sv:10:5
										localparam BLOCK_SIZE = 1;
										// Trace: src/VX_fpu_unit.sv:11:5
										localparam NUM_LANES = 4;
										// Trace: src/VX_fpu_unit.sv:12:5
										localparam PID_BITS = 0;
										// Trace: src/VX_fpu_unit.sv:13:5
										localparam PID_WIDTH = 1;
										// Trace: src/VX_fpu_unit.sv:14:5
										localparam TAG_WIDTH = 1;
										// Trace: src/VX_fpu_unit.sv:15:5
										localparam PARTIAL_BW = 1'd0;
										// Trace: src/VX_fpu_unit.sv:16:5
										// expanded interface instance: per_block_execute_if
										localparam _param_E2592_NUM_LANES = NUM_LANES;
										genvar _arr_E2592;
										for (_arr_E2592 = 0; _arr_E2592 <= 0; _arr_E2592 = _arr_E2592 + 1) begin : per_block_execute_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_execute_if.sv:2:15
											localparam NUM_LANES = _param_E2592_NUM_LANES;
											// Trace: src/VX_execute_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_execute_if.sv:5:5
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_execute_if.sv:22:5
											wire valid;
											// Trace: src/VX_execute_if.sv:23:5
											wire [474:0] data;
											// Trace: src/VX_execute_if.sv:24:5
											wire ready;
											// Trace: src/VX_execute_if.sv:25:5
											// Trace: src/VX_execute_if.sv:30:5
										end
										// Trace: src/VX_fpu_unit.sv:19:5
										// expanded module instance: dispatch_unit
										localparam _bbase_2E16E_dispatch_if = 3;
										localparam _bbase_2E16E_execute_if = 0;
										localparam _param_2E16E_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_2E16E_NUM_LANES = NUM_LANES;
										localparam _param_2E16E_OUT_BUF = (PARTIAL_BW ? 3 : 0);
										if (1) begin : dispatch_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_dispatch_unit.sv:2:15
											localparam BLOCK_SIZE = _param_2E16E_BLOCK_SIZE;
											// Trace: src/VX_dispatch_unit.sv:3:15
											localparam NUM_LANES = _param_2E16E_NUM_LANES;
											// Trace: src/VX_dispatch_unit.sv:4:15
											localparam OUT_BUF = _param_2E16E_OUT_BUF;
											// Trace: src/VX_dispatch_unit.sv:5:15
											localparam MAX_FANOUT = 8;
											// Trace: src/VX_dispatch_unit.sv:7:5
											wire clk;
											// Trace: src/VX_dispatch_unit.sv:8:5
											wire reset;
											// Trace: src/VX_dispatch_unit.sv:9:5
											localparam _mbase_dispatch_if = 3;
											// Trace: src/VX_dispatch_unit.sv:10:5
											localparam _mbase_execute_if = 0;
											// Trace: src/VX_dispatch_unit.sv:12:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:13:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_dispatch_unit.sv:14:5
											localparam PID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:15:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:16:5
											localparam BATCH_COUNT = 1;
											// Trace: src/VX_dispatch_unit.sv:17:5
											localparam BATCH_COUNT_W = 1;
											// Trace: src/VX_dispatch_unit.sv:18:5
											localparam ISSUE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:19:5
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											localparam VX_gpu_pkg_ISSUE_WIS = 2;
											localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											localparam IN_DATAW = 472;
											// Trace: src/VX_dispatch_unit.sv:20:5
											localparam OUT_DATAW = 475;
											// Trace: src/VX_dispatch_unit.sv:21:5
											localparam FANOUT_ENABLE = 1'd0;
											// Trace: src/VX_dispatch_unit.sv:22:5
											localparam DATA_TMASK_OFF = 465;
											// Trace: src/VX_dispatch_unit.sv:23:5
											localparam DATA_REGS_OFF = 0;
											// Trace: src/VX_dispatch_unit.sv:24:5
											wire [0:0] dispatch_valid;
											// Trace: src/VX_dispatch_unit.sv:25:5
											wire [471:0] dispatch_data;
											// Trace: src/VX_dispatch_unit.sv:26:5
											wire [0:0] dispatch_ready;
											// Trace: src/VX_dispatch_unit.sv:27:5
											genvar _gv_i_96;
											for (_gv_i_96 = 0; _gv_i_96 < 1; _gv_i_96 = _gv_i_96 + 1) begin : g_dispatch_data
												localparam i = _gv_i_96;
												// Trace: src/VX_dispatch_unit.sv:28:9
												assign dispatch_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].valid;
												// Trace: src/VX_dispatch_unit.sv:29:9
												assign dispatch_data[i * 472+:472] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].data;
												// Trace: src/VX_dispatch_unit.sv:30:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].ready = dispatch_ready[i];
											end
											// Trace: src/VX_dispatch_unit.sv:32:5
											wire [0:0] block_ready;
											// Trace: src/VX_dispatch_unit.sv:33:5
											wire [3:0] block_tmask;
											// Trace: src/VX_dispatch_unit.sv:34:5
											wire [383:0] block_regs;
											// Trace: src/VX_dispatch_unit.sv:35:5
											wire [0:0] block_pid;
											// Trace: src/VX_dispatch_unit.sv:36:5
											wire [0:0] block_sop;
											// Trace: src/VX_dispatch_unit.sv:37:5
											wire [0:0] block_eop;
											// Trace: src/VX_dispatch_unit.sv:38:5
											wire [0:0] block_done;
											// Trace: src/VX_dispatch_unit.sv:39:5
											wire batch_done = &block_done;
											// Trace: src/VX_dispatch_unit.sv:40:5
											wire [0:0] batch_idx;
											// Trace: src/VX_dispatch_unit.sv:41:5
											if (1) begin : g_batch_idx_0
												// Trace: src/VX_dispatch_unit.sv:67:9
												assign batch_idx = 0;
											end
											// Trace: src/VX_dispatch_unit.sv:69:5
											wire [0:0] issue_indices;
											// Trace: src/VX_dispatch_unit.sv:70:5
											genvar _gv_block_idx_2;
											for (_gv_block_idx_2 = 0; _gv_block_idx_2 < BLOCK_SIZE; _gv_block_idx_2 = _gv_block_idx_2 + 1) begin : g_issue_indices
												localparam block_idx = _gv_block_idx_2;
												// Trace: src/VX_dispatch_unit.sv:71:9
												assign issue_indices[block_idx+:1] = sv2v_cast_1(batch_idx * BLOCK_SIZE) + sv2v_cast_1_signed(block_idx);
											end
											// Trace: src/VX_dispatch_unit.sv:73:5
											genvar _gv_block_idx_3;
											localparam VX_gpu_pkg_ISSUE_ISW = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											function [1:0] VX_gpu_pkg_wis_to_wid;
												// Trace: src/VX_gpu_pkg.sv:151:9
												input reg [1:0] wis;
												// Trace: src/VX_gpu_pkg.sv:152:9
												input reg [0:0] isw;
												// Trace: src/VX_gpu_pkg.sv:154:9
												begin
													// Trace: src/VX_gpu_pkg.sv:157:13
													VX_gpu_pkg_wis_to_wid = wis;
												end
											endfunction
											for (_gv_block_idx_3 = 0; _gv_block_idx_3 < BLOCK_SIZE; _gv_block_idx_3 = _gv_block_idx_3 + 1) begin : g_blocks
												localparam block_idx = _gv_block_idx_3;
												// Trace: src/VX_dispatch_unit.sv:74:9
												wire [0:0] issue_idx = issue_indices[block_idx+:1];
												// Trace: src/VX_dispatch_unit.sv:75:9
												wire valid_p;
												wire ready_p;
												if (1) begin : g_full_threads
													// Trace: src/VX_dispatch_unit.sv:168:13
													assign valid_p = dispatch_valid[issue_idx];
													// Trace: src/VX_dispatch_unit.sv:169:13
													assign block_tmask[block_idx * 4+:4] = dispatch_data[(issue_idx * 472) + DATA_TMASK_OFF+:4];
													// Trace: src/VX_dispatch_unit.sv:170:13
													assign block_regs[32 * ((block_idx * 3) * 4)+:128] = dispatch_data[(issue_idx * 472) + 256+:128];
													// Trace: src/VX_dispatch_unit.sv:171:13
													assign block_regs[32 * (((block_idx * 3) + 1) * 4)+:128] = dispatch_data[(issue_idx * 472) + 128+:128];
													// Trace: src/VX_dispatch_unit.sv:172:13
													assign block_regs[32 * (((block_idx * 3) + 2) * 4)+:128] = dispatch_data[issue_idx * 472+:128];
													// Trace: src/VX_dispatch_unit.sv:173:13
													assign block_pid[block_idx+:1] = 1'sb0;
													// Trace: src/VX_dispatch_unit.sv:174:13
													assign block_sop[block_idx] = 1'b1;
													// Trace: src/VX_dispatch_unit.sv:175:13
													assign block_eop[block_idx] = 1'b1;
													// Trace: src/VX_dispatch_unit.sv:176:13
													assign block_ready[block_idx] = ready_p;
													// Trace: src/VX_dispatch_unit.sv:177:13
													assign block_done[block_idx] = ready_p || ~valid_p;
												end
												// Trace: src/VX_dispatch_unit.sv:179:9
												wire [0:0] isw;
												if (1) begin : g_isw
													// Trace: src/VX_dispatch_unit.sv:187:13
													assign isw = block_idx;
												end
												// Trace: src/VX_dispatch_unit.sv:189:9
												wire [1:0] block_wid = VX_gpu_pkg_wis_to_wid(dispatch_data[(issue_idx * 472) + 469+:VX_gpu_pkg_ISSUE_WIS_W], isw);
												// Trace: src/VX_dispatch_unit.sv:190:9
												wire [474:0] execute_data;
												reg [474:0] execute_data_w;
												// Trace: src/VX_dispatch_unit.sv:191:9
												VX_elastic_buffer #(
													.DATAW(OUT_DATAW),
													.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
													.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
												) buf_out(
													.clk(clk),
													.reset(reset),
													.valid_in(valid_p),
													.ready_in(ready_p),
													.data_in({dispatch_data[(issue_idx * 472) + 471-:1], block_wid, block_tmask[block_idx * 4+:4], dispatch_data[(issue_idx * 472) + 464-:81], block_regs[32 * ((block_idx * 3) * 4)+:128], block_regs[32 * (((block_idx * 3) + 1) * 4)+:128], block_regs[32 * (((block_idx * 3) + 2) * 4)+:128], block_pid[block_idx+:1], block_sop[block_idx], block_eop[block_idx]}),
													.data_out(execute_data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_unit.per_block_execute_if[block_idx + _mbase_execute_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_unit.per_block_execute_if[block_idx + _mbase_execute_if].ready)
												);
												if (1) begin : g_execute_data_w_full
													// Trace: src/VX_dispatch_unit.sv:218:13
													always @(*) begin
														// Trace: src/VX_dispatch_unit.sv:219:17
														execute_data_w = execute_data;
														// Trace: src/VX_dispatch_unit.sv:220:17
														execute_data_w[2:0] = 3'b011;
													end
												end
												// Trace: src/VX_dispatch_unit.sv:223:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_unit.per_block_execute_if[block_idx + _mbase_execute_if].data = execute_data_w;
											end
											// Trace: src/VX_dispatch_unit.sv:225:5
											reg [0:0] ready_in;
											// Trace: src/VX_dispatch_unit.sv:226:5
											always @(*) begin
												// Trace: src/VX_dispatch_unit.sv:227:9
												ready_in = 0;
												// Trace: src/VX_dispatch_unit.sv:228:9
												begin : sv2v_autoblock_15
													// Trace: src/VX_dispatch_unit.sv:228:14
													integer block_idx;
													// Trace: src/VX_dispatch_unit.sv:228:14
													for (block_idx = 0; block_idx < BLOCK_SIZE; block_idx = block_idx + 1)
														begin
															// Trace: src/VX_dispatch_unit.sv:229:13
															ready_in[issue_indices[block_idx+:1]] = block_ready[block_idx] && block_eop[block_idx];
														end
												end
											end
											// Trace: src/VX_dispatch_unit.sv:232:5
											assign dispatch_ready = ready_in;
										end
										assign dispatch_unit.clk = clk;
										assign dispatch_unit.reset = reset;
										// Trace: src/VX_fpu_unit.sv:29:5
										// expanded interface instance: per_block_commit_if
										localparam _param_98792_NUM_LANES = NUM_LANES;
										genvar _arr_98792;
										for (_arr_98792 = 0; _arr_98792 <= 0; _arr_98792 = _arr_98792 + 1) begin : per_block_commit_if
											// Trace: src/VX_commit_if.sv:2:15
											localparam NUM_LANES = _param_98792_NUM_LANES;
											// Trace: src/VX_commit_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_commit_if.sv:5:5
											// removed localparam type data_t
											// Trace: src/VX_commit_if.sv:17:5
											wire valid;
											// Trace: src/VX_commit_if.sv:18:5
											wire [175:0] data;
											// Trace: src/VX_commit_if.sv:19:5
											wire ready;
											// Trace: src/VX_commit_if.sv:20:5
											// Trace: src/VX_commit_if.sv:25:5
										end
										// Trace: src/VX_fpu_unit.sv:32:5
										genvar _gv_block_idx_4;
										// removed localparam type VX_fpu_pkg_fflags_t
										for (_gv_block_idx_4 = 0; _gv_block_idx_4 < BLOCK_SIZE; _gv_block_idx_4 = _gv_block_idx_4 + 1) begin : g_fpus
											localparam block_idx = _gv_block_idx_4;
											// Trace: src/VX_fpu_unit.sv:33:9
											wire fpu_req_valid;
											wire fpu_req_ready;
											// Trace: src/VX_fpu_unit.sv:34:9
											wire fpu_rsp_valid;
											wire fpu_rsp_ready;
											// Trace: src/VX_fpu_unit.sv:35:9
											wire [127:0] fpu_rsp_result;
											// Trace: src/VX_fpu_unit.sv:36:9
											wire [4:0] fpu_rsp_fflags;
											// Trace: src/VX_fpu_unit.sv:37:9
											wire fpu_rsp_has_fflags;
											// Trace: src/VX_fpu_unit.sv:38:9
											wire [0:0] fpu_rsp_uuid;
											// Trace: src/VX_fpu_unit.sv:39:9
											wire [1:0] fpu_rsp_wid;
											// Trace: src/VX_fpu_unit.sv:40:9
											wire [3:0] fpu_rsp_tmask;
											// Trace: src/VX_fpu_unit.sv:41:9
											wire [30:0] fpu_rsp_PC;
											// Trace: src/VX_fpu_unit.sv:42:9
											wire [5:0] fpu_rsp_rd;
											// Trace: src/VX_fpu_unit.sv:43:9
											wire [0:0] fpu_rsp_pid;
											wire [0:0] fpu_rsp_pid_u;
											// Trace: src/VX_fpu_unit.sv:44:9
											wire fpu_rsp_sop;
											wire fpu_rsp_sop_u;
											// Trace: src/VX_fpu_unit.sv:45:9
											wire fpu_rsp_eop;
											wire fpu_rsp_eop_u;
											// Trace: src/VX_fpu_unit.sv:46:9
											wire [0:0] fpu_req_tag;
											wire [0:0] fpu_rsp_tag;
											// Trace: src/VX_fpu_unit.sv:47:9
											wire mdata_full;
											// Trace: src/VX_fpu_unit.sv:48:9
											wire [1:0] fpu_fmt = per_block_execute_if[block_idx].data[397-:2];
											// Trace: src/VX_fpu_unit.sv:49:9
											wire [2:0] fpu_frm = per_block_execute_if[block_idx].data[400-:3];
											// Trace: src/VX_fpu_unit.sv:50:9
											wire execute_fire = per_block_execute_if[block_idx].valid && per_block_execute_if[block_idx].ready;
											// Trace: src/VX_fpu_unit.sv:51:9
											wire fpu_rsp_fire = fpu_rsp_valid && fpu_rsp_ready;
											// Trace: src/VX_fpu_unit.sv:52:9
											VX_index_buffer #(
												.DATAW(47),
												.SIZE(2)
											) tag_store(
												.clk(clk),
												.reset(reset),
												.acquire_en(execute_fire),
												.write_addr(fpu_req_tag),
												.write_data({per_block_execute_if[block_idx].data[474], per_block_execute_if[block_idx].data[473-:2], per_block_execute_if[block_idx].data[471-:4], per_block_execute_if[block_idx].data[467-:31], per_block_execute_if[block_idx].data[394-:6], per_block_execute_if[block_idx].data[2], per_block_execute_if[block_idx].data[1], per_block_execute_if[block_idx].data[0]}),
												.read_data({fpu_rsp_uuid, fpu_rsp_wid, fpu_rsp_tmask, fpu_rsp_PC, fpu_rsp_rd, fpu_rsp_pid_u, fpu_rsp_sop_u, fpu_rsp_eop_u}),
												.read_addr(fpu_rsp_tag),
												.release_en(fpu_rsp_fire),
												.full(mdata_full),
												.empty()
											);
											if (1) begin : g_no_fpu_rsp_pid
												// Trace: src/VX_fpu_unit.sv:72:13
												assign fpu_rsp_pid = 0;
												// Trace: src/VX_fpu_unit.sv:73:13
												assign fpu_rsp_sop = 1;
												// Trace: src/VX_fpu_unit.sv:74:13
												assign fpu_rsp_eop = 1;
											end
											// Trace: src/VX_fpu_unit.sv:76:9
											wire [2:0] fpu_req_frm;
											if (1) begin : genblk2
												// Trace: src/VX_fpu_unit.sv:85:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[block_idx + _mbase_fpu_csr_if].read_wid = per_block_execute_if[block_idx].data[473-:2];
											end
											// Trace: src/VX_fpu_unit.sv:88:9
											assign fpu_req_frm = ((per_block_execute_if[block_idx].data[436-:4] != 4'b1110) && (fpu_frm == 3'b111) ? Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[block_idx + _mbase_fpu_csr_if].read_frm : fpu_frm);
											// Trace: src/VX_fpu_unit.sv:90:9
											assign fpu_req_valid = per_block_execute_if[block_idx].valid && ~mdata_full;
											// Trace: src/VX_fpu_unit.sv:91:9
											assign per_block_execute_if[block_idx].ready = fpu_req_ready && ~mdata_full;
											// Trace: src/VX_fpu_unit.sv:92:9
											VX_fpu_fpnew #(
												.NUM_LANES(NUM_LANES),
												.TAG_WIDTH(TAG_WIDTH),
												.OUT_BUF((PARTIAL_BW ? 1 : 3))
											) fpu_fpnew(
												.clk(clk),
												.reset(reset),
												.valid_in(fpu_req_valid),
												.mask_in(per_block_execute_if[block_idx].data[471-:4]),
												.op_type(per_block_execute_if[block_idx].data[436-:4]),
												.fmt(fpu_fmt),
												.frm(fpu_req_frm),
												.dataa(per_block_execute_if[block_idx].data[386-:128]),
												.datab(per_block_execute_if[block_idx].data[258-:128]),
												.datac(per_block_execute_if[block_idx].data[130-:128]),
												.tag_in(fpu_req_tag),
												.ready_in(fpu_req_ready),
												.valid_out(fpu_rsp_valid),
												.result(fpu_rsp_result),
												.has_fflags(fpu_rsp_has_fflags),
												.fflags(fpu_rsp_fflags),
												.tag_out(fpu_rsp_tag),
												.ready_out(fpu_rsp_ready)
											);
											// Trace: src/VX_fpu_unit.sv:116:9
											wire [4:0] fpu_rsp_fflags_q;
											if (1) begin : g_no_pid
												// Trace: src/VX_fpu_unit.sv:128:13
												assign fpu_rsp_fflags_q = fpu_rsp_fflags;
											end
											// Trace: src/VX_fpu_unit.sv:130:9
											// expanded interface instance: fpu_csr_tmp_if
											if (1) begin : fpu_csr_tmp_if
												// removed import VX_fpu_pkg::*;
												// Trace: src/VX_fpu_csr_if.sv:2:5
												wire write_enable;
												// Trace: src/VX_fpu_csr_if.sv:3:5
												wire [1:0] write_wid;
												// Trace: src/VX_fpu_csr_if.sv:4:5
												// removed localparam type VX_fpu_pkg_fflags_t
												wire [4:0] write_fflags;
												// Trace: src/VX_fpu_csr_if.sv:5:5
												wire [1:0] read_wid;
												// Trace: src/VX_fpu_csr_if.sv:6:5
												wire [2:0] read_frm;
												// Trace: src/VX_fpu_csr_if.sv:7:5
												// Trace: src/VX_fpu_csr_if.sv:14:5
											end
											// Trace: src/VX_fpu_unit.sv:131:9
											assign fpu_csr_tmp_if.write_enable = (fpu_rsp_fire && fpu_rsp_eop) && fpu_rsp_has_fflags;
											if (1) begin : genblk4
												// Trace: src/VX_fpu_unit.sv:140:9
												assign fpu_csr_tmp_if.write_wid = fpu_rsp_wid;
											end
											// Trace: src/VX_fpu_unit.sv:143:9
											assign fpu_csr_tmp_if.write_fflags = fpu_rsp_fflags_q;
											// Trace: src/VX_fpu_unit.sv:144:10
											VX_pipe_register #(
												.DATAW(8),
												.RESETW(1)
											) fpu_csr_reg(
												.clk(clk),
												.reset(reset),
												.enable(1'b1),
												.data_in({fpu_csr_tmp_if.write_enable, fpu_csr_tmp_if.write_wid, fpu_csr_tmp_if.write_fflags}),
												.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[block_idx + _mbase_fpu_csr_if].write_enable, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[block_idx + _mbase_fpu_csr_if].write_wid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[block_idx + _mbase_fpu_csr_if].write_fflags})
											);
											// Trace: src/VX_fpu_unit.sv:154:9
											VX_elastic_buffer #(
												.DATAW(175),
												.SIZE(0)
											) rsp_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(fpu_rsp_valid),
												.ready_in(fpu_rsp_ready),
												.data_in({fpu_rsp_uuid, fpu_rsp_wid, fpu_rsp_tmask, fpu_rsp_PC, fpu_rsp_rd, fpu_rsp_result, fpu_rsp_pid, fpu_rsp_sop, fpu_rsp_eop}),
												.data_out({per_block_commit_if[block_idx].data[175], per_block_commit_if[block_idx].data[174-:2], per_block_commit_if[block_idx].data[172-:4], per_block_commit_if[block_idx].data[168-:31], per_block_commit_if[block_idx].data[136-:6], per_block_commit_if[block_idx].data[130-:128], per_block_commit_if[block_idx].data[2], per_block_commit_if[block_idx].data[1], per_block_commit_if[block_idx].data[0]}),
												.valid_out(per_block_commit_if[block_idx].valid),
												.ready_out(per_block_commit_if[block_idx].ready)
											);
											// Trace: src/VX_fpu_unit.sv:167:9
											assign per_block_commit_if[block_idx].data[137] = 1'b1;
										end
										// Trace: src/VX_fpu_unit.sv:169:5
										// expanded module instance: gather_unit
										localparam _bbase_8E516_commit_in_if = 0;
										localparam _bbase_8E516_commit_out_if = 3;
										localparam _param_8E516_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_8E516_NUM_LANES = NUM_LANES;
										localparam _param_8E516_OUT_BUF = (PARTIAL_BW ? 3 : 0);
										if (1) begin : gather_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_gather_unit.sv:2:15
											localparam BLOCK_SIZE = _param_8E516_BLOCK_SIZE;
											// Trace: src/VX_gather_unit.sv:3:15
											localparam NUM_LANES = _param_8E516_NUM_LANES;
											// Trace: src/VX_gather_unit.sv:4:15
											localparam OUT_BUF = _param_8E516_OUT_BUF;
											// Trace: src/VX_gather_unit.sv:6:5
											wire clk;
											// Trace: src/VX_gather_unit.sv:7:5
											wire reset;
											// Trace: src/VX_gather_unit.sv:8:5
											localparam _mbase_commit_in_if = 0;
											// Trace: src/VX_gather_unit.sv:9:5
											localparam _mbase_commit_out_if = 3;
											// Trace: src/VX_gather_unit.sv:11:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_gather_unit.sv:12:5
											localparam PID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:13:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:14:5
											localparam DATAW = 176;
											// Trace: src/VX_gather_unit.sv:15:5
											localparam DATA_WIS_OFF = 173;
											// Trace: src/VX_gather_unit.sv:16:5
											wire [0:0] commit_in_valid;
											// Trace: src/VX_gather_unit.sv:17:5
											wire [175:0] commit_in_data;
											// Trace: src/VX_gather_unit.sv:18:5
											wire [0:0] commit_in_ready;
											// Trace: src/VX_gather_unit.sv:19:5
											localparam VX_gpu_pkg_ISSUE_ISW = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											wire [0:0] commit_in_isw;
											// Trace: src/VX_gather_unit.sv:20:5
											genvar _gv_i_208;
											for (_gv_i_208 = 0; _gv_i_208 < BLOCK_SIZE; _gv_i_208 = _gv_i_208 + 1) begin : g_commit_in
												localparam i = _gv_i_208;
												// Trace: src/VX_gather_unit.sv:21:9
												assign commit_in_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_unit.per_block_commit_if[i + _mbase_commit_in_if].valid;
												// Trace: src/VX_gather_unit.sv:22:9
												assign commit_in_data[i * 176+:176] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_unit.per_block_commit_if[i + _mbase_commit_in_if].data;
												// Trace: src/VX_gather_unit.sv:23:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_unit.per_block_commit_if[i + _mbase_commit_in_if].ready = commit_in_ready[i];
												if (1) begin : g_commit_in_isw_full
													// Trace: src/VX_gather_unit.sv:31:13
													assign commit_in_isw[i+:1] = sv2v_cast_1_signed(i);
												end
											end
											// Trace: src/VX_gather_unit.sv:34:5
											reg [0:0] commit_out_valid;
											// Trace: src/VX_gather_unit.sv:35:5
											reg [175:0] commit_out_data;
											// Trace: src/VX_gather_unit.sv:36:5
											wire [0:0] commit_out_ready;
											// Trace: src/VX_gather_unit.sv:37:5
											always @(*) begin
												// Trace: src/VX_gather_unit.sv:38:9
												commit_out_valid = 1'sb0;
												// Trace: src/VX_gather_unit.sv:39:9
												begin : sv2v_autoblock_16
													// Trace: src/VX_gather_unit.sv:39:14
													integer i;
													// Trace: src/VX_gather_unit.sv:39:14
													for (i = 0; i < 1; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:40:13
															commit_out_data[i * 176+:176] = 1'sbx;
														end
												end
												begin : sv2v_autoblock_17
													// Trace: src/VX_gather_unit.sv:42:14
													integer i;
													// Trace: src/VX_gather_unit.sv:42:14
													for (i = 0; i < BLOCK_SIZE; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:43:13
															commit_out_valid[commit_in_isw[i+:1]] = commit_in_valid[i];
															// Trace: src/VX_gather_unit.sv:44:13
															commit_out_data[commit_in_isw[i+:1] * 176+:176] = commit_in_data[i * 176+:176];
														end
												end
											end
											// Trace: src/VX_gather_unit.sv:47:5
											genvar _gv_i_209;
											for (_gv_i_209 = 0; _gv_i_209 < BLOCK_SIZE; _gv_i_209 = _gv_i_209 + 1) begin : g_commit_in_ready
												localparam i = _gv_i_209;
												// Trace: src/VX_gather_unit.sv:48:9
												assign commit_in_ready[i] = commit_out_ready[commit_in_isw[i+:1]];
											end
											// Trace: src/VX_gather_unit.sv:50:5
											genvar _gv_i_210;
											for (_gv_i_210 = 0; _gv_i_210 < 1; _gv_i_210 = _gv_i_210 + 1) begin : g_out_bufs
												localparam i = _gv_i_210;
												// Trace: src/VX_gather_unit.sv:51:9
												// expanded interface instance: commit_tmp_if
												localparam _param_C9958_NUM_LANES = NUM_LANES;
												if (1) begin : commit_tmp_if
													// Trace: src/VX_commit_if.sv:2:15
													localparam NUM_LANES = _param_C9958_NUM_LANES;
													// Trace: src/VX_commit_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_commit_if.sv:5:5
													// removed localparam type data_t
													// Trace: src/VX_commit_if.sv:17:5
													wire valid;
													// Trace: src/VX_commit_if.sv:18:5
													wire [175:0] data;
													// Trace: src/VX_commit_if.sv:19:5
													wire ready;
													// Trace: src/VX_commit_if.sv:20:5
													// Trace: src/VX_commit_if.sv:25:5
												end
												// Trace: src/VX_gather_unit.sv:54:9
												VX_elastic_buffer #(
													.DATAW(DATAW),
													.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
													.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
												) out_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(commit_out_valid[i]),
													.ready_in(commit_out_ready[i]),
													.data_in(commit_out_data[i * 176+:176]),
													.data_out(commit_tmp_if.data),
													.valid_out(commit_tmp_if.valid),
													.ready_out(commit_tmp_if.ready)
												);
												// Trace: src/VX_gather_unit.sv:68:9
												wire [3:0] commit_tmask_w;
												// Trace: src/VX_gather_unit.sv:69:9
												wire [127:0] commit_data_w;
												if (1) begin : g_commit_data_no_pid
													// Trace: src/VX_gather_unit.sv:80:13
													assign commit_tmask_w = commit_tmp_if.data[172-:4];
													// Trace: src/VX_gather_unit.sv:81:13
													assign commit_data_w = commit_tmp_if.data[130-:128];
												end
												// Trace: src/VX_gather_unit.sv:83:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].valid = commit_tmp_if.valid;
												// Trace: src/VX_gather_unit.sv:84:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].data = {commit_tmp_if.data[175], commit_tmp_if.data[174-:2], commit_tmask_w, commit_tmp_if.data[168-:31], commit_tmp_if.data[137], commit_tmp_if.data[136-:6], commit_data_w, 1'b0, commit_tmp_if.data[1], commit_tmp_if.data[0]};
												// Trace: src/VX_gather_unit.sv:96:9
												assign commit_tmp_if.ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].ready;
											end
										end
										assign gather_unit.clk = clk;
										assign gather_unit.reset = reset;
									end
									assign fpu_unit.clk = clk;
									assign fpu_unit.reset = reset;
									// Trace: src/VX_execute.sv:45:5
									// expanded module instance: sfu_unit
									localparam _bbase_6660E_dispatch_if = 2;
									localparam _bbase_6660E_commit_if = 2;
									localparam _bbase_6660E_fpu_csr_if = 0;
									localparam _param_6660E_INSTANCE_ID = "";
									localparam _param_6660E_CORE_ID = CORE_ID;
									if (1) begin : sfu_unit
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_sfu_unit.sv:2:16
										localparam INSTANCE_ID = _param_6660E_INSTANCE_ID;
										// Trace: src/VX_sfu_unit.sv:3:15
										localparam CORE_ID = _param_6660E_CORE_ID;
										// Trace: src/VX_sfu_unit.sv:5:5
										wire clk;
										// Trace: src/VX_sfu_unit.sv:6:5
										wire reset;
										// Trace: src/VX_sfu_unit.sv:7:5
										// removed localparam type VX_gpu_pkg_base_dcrs_t
										wire [71:0] base_dcrs;
										// Trace: src/VX_sfu_unit.sv:8:5
										localparam _mbase_dispatch_if = 2;
										// Trace: src/VX_sfu_unit.sv:9:5
										localparam _mbase_fpu_csr_if = 0;
										// Trace: src/VX_sfu_unit.sv:10:5
										// removed modport instance commit_csr_if
										// Trace: src/VX_sfu_unit.sv:11:5
										// removed modport instance sched_csr_if
										// Trace: src/VX_sfu_unit.sv:12:5
										localparam _mbase_commit_if = 2;
										// Trace: src/VX_sfu_unit.sv:13:5
										// removed modport instance warp_ctl_if
										// Trace: src/VX_sfu_unit.sv:15:5
										localparam BLOCK_SIZE = 1;
										// Trace: src/VX_sfu_unit.sv:16:5
										localparam NUM_LANES = 4;
										// Trace: src/VX_sfu_unit.sv:17:5
										localparam PE_COUNT = 2;
										// Trace: src/VX_sfu_unit.sv:18:5
										localparam PE_SEL_BITS = 1;
										// Trace: src/VX_sfu_unit.sv:19:5
										localparam PE_IDX_WCTL = 0;
										// Trace: src/VX_sfu_unit.sv:20:5
										localparam PE_IDX_CSRS = 1;
										// Trace: src/VX_sfu_unit.sv:21:5
										// expanded interface instance: per_block_execute_if
										localparam _param_E2592_NUM_LANES = NUM_LANES;
										genvar _arr_E2592;
										for (_arr_E2592 = 0; _arr_E2592 <= 0; _arr_E2592 = _arr_E2592 + 1) begin : per_block_execute_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_execute_if.sv:2:15
											localparam NUM_LANES = _param_E2592_NUM_LANES;
											// Trace: src/VX_execute_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_execute_if.sv:5:5
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_execute_if.sv:22:5
											wire valid;
											// Trace: src/VX_execute_if.sv:23:5
											wire [474:0] data;
											// Trace: src/VX_execute_if.sv:24:5
											wire ready;
											// Trace: src/VX_execute_if.sv:25:5
											// Trace: src/VX_execute_if.sv:30:5
										end
										// Trace: src/VX_sfu_unit.sv:24:5
										// expanded interface instance: per_block_commit_if
										localparam _param_98792_NUM_LANES = NUM_LANES;
										genvar _arr_98792;
										for (_arr_98792 = 0; _arr_98792 <= 0; _arr_98792 = _arr_98792 + 1) begin : per_block_commit_if
											// Trace: src/VX_commit_if.sv:2:15
											localparam NUM_LANES = _param_98792_NUM_LANES;
											// Trace: src/VX_commit_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_commit_if.sv:5:5
											// removed localparam type data_t
											// Trace: src/VX_commit_if.sv:17:5
											wire valid;
											// Trace: src/VX_commit_if.sv:18:5
											wire [175:0] data;
											// Trace: src/VX_commit_if.sv:19:5
											wire ready;
											// Trace: src/VX_commit_if.sv:20:5
											// Trace: src/VX_commit_if.sv:25:5
										end
										// Trace: src/VX_sfu_unit.sv:27:5
										// expanded module instance: dispatch_unit
										localparam _bbase_2E16E_dispatch_if = 2;
										localparam _bbase_2E16E_execute_if = 0;
										localparam _param_2E16E_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_2E16E_NUM_LANES = NUM_LANES;
										localparam _param_2E16E_OUT_BUF = 3;
										if (1) begin : dispatch_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_dispatch_unit.sv:2:15
											localparam BLOCK_SIZE = _param_2E16E_BLOCK_SIZE;
											// Trace: src/VX_dispatch_unit.sv:3:15
											localparam NUM_LANES = _param_2E16E_NUM_LANES;
											// Trace: src/VX_dispatch_unit.sv:4:15
											localparam OUT_BUF = _param_2E16E_OUT_BUF;
											// Trace: src/VX_dispatch_unit.sv:5:15
											localparam MAX_FANOUT = 8;
											// Trace: src/VX_dispatch_unit.sv:7:5
											wire clk;
											// Trace: src/VX_dispatch_unit.sv:8:5
											wire reset;
											// Trace: src/VX_dispatch_unit.sv:9:5
											localparam _mbase_dispatch_if = 2;
											// Trace: src/VX_dispatch_unit.sv:10:5
											localparam _mbase_execute_if = 0;
											// Trace: src/VX_dispatch_unit.sv:12:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:13:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_dispatch_unit.sv:14:5
											localparam PID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:15:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:16:5
											localparam BATCH_COUNT = 1;
											// Trace: src/VX_dispatch_unit.sv:17:5
											localparam BATCH_COUNT_W = 1;
											// Trace: src/VX_dispatch_unit.sv:18:5
											localparam ISSUE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:19:5
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											localparam VX_gpu_pkg_ISSUE_WIS = 2;
											localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											localparam IN_DATAW = 472;
											// Trace: src/VX_dispatch_unit.sv:20:5
											localparam OUT_DATAW = 475;
											// Trace: src/VX_dispatch_unit.sv:21:5
											localparam FANOUT_ENABLE = 1'd0;
											// Trace: src/VX_dispatch_unit.sv:22:5
											localparam DATA_TMASK_OFF = 465;
											// Trace: src/VX_dispatch_unit.sv:23:5
											localparam DATA_REGS_OFF = 0;
											// Trace: src/VX_dispatch_unit.sv:24:5
											wire [0:0] dispatch_valid;
											// Trace: src/VX_dispatch_unit.sv:25:5
											wire [471:0] dispatch_data;
											// Trace: src/VX_dispatch_unit.sv:26:5
											wire [0:0] dispatch_ready;
											// Trace: src/VX_dispatch_unit.sv:27:5
											genvar _gv_i_96;
											for (_gv_i_96 = 0; _gv_i_96 < 1; _gv_i_96 = _gv_i_96 + 1) begin : g_dispatch_data
												localparam i = _gv_i_96;
												// Trace: src/VX_dispatch_unit.sv:28:9
												assign dispatch_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].valid;
												// Trace: src/VX_dispatch_unit.sv:29:9
												assign dispatch_data[i * 472+:472] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].data;
												// Trace: src/VX_dispatch_unit.sv:30:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].ready = dispatch_ready[i];
											end
											// Trace: src/VX_dispatch_unit.sv:32:5
											wire [0:0] block_ready;
											// Trace: src/VX_dispatch_unit.sv:33:5
											wire [3:0] block_tmask;
											// Trace: src/VX_dispatch_unit.sv:34:5
											wire [383:0] block_regs;
											// Trace: src/VX_dispatch_unit.sv:35:5
											wire [0:0] block_pid;
											// Trace: src/VX_dispatch_unit.sv:36:5
											wire [0:0] block_sop;
											// Trace: src/VX_dispatch_unit.sv:37:5
											wire [0:0] block_eop;
											// Trace: src/VX_dispatch_unit.sv:38:5
											wire [0:0] block_done;
											// Trace: src/VX_dispatch_unit.sv:39:5
											wire batch_done = &block_done;
											// Trace: src/VX_dispatch_unit.sv:40:5
											wire [0:0] batch_idx;
											// Trace: src/VX_dispatch_unit.sv:41:5
											if (1) begin : g_batch_idx_0
												// Trace: src/VX_dispatch_unit.sv:67:9
												assign batch_idx = 0;
											end
											// Trace: src/VX_dispatch_unit.sv:69:5
											wire [0:0] issue_indices;
											// Trace: src/VX_dispatch_unit.sv:70:5
											genvar _gv_block_idx_2;
											for (_gv_block_idx_2 = 0; _gv_block_idx_2 < BLOCK_SIZE; _gv_block_idx_2 = _gv_block_idx_2 + 1) begin : g_issue_indices
												localparam block_idx = _gv_block_idx_2;
												// Trace: src/VX_dispatch_unit.sv:71:9
												assign issue_indices[block_idx+:1] = sv2v_cast_1(batch_idx * BLOCK_SIZE) + sv2v_cast_1_signed(block_idx);
											end
											// Trace: src/VX_dispatch_unit.sv:73:5
											genvar _gv_block_idx_3;
											localparam VX_gpu_pkg_ISSUE_ISW = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											function [1:0] VX_gpu_pkg_wis_to_wid;
												// Trace: src/VX_gpu_pkg.sv:151:9
												input reg [1:0] wis;
												// Trace: src/VX_gpu_pkg.sv:152:9
												input reg [0:0] isw;
												// Trace: src/VX_gpu_pkg.sv:154:9
												begin
													// Trace: src/VX_gpu_pkg.sv:157:13
													VX_gpu_pkg_wis_to_wid = wis;
												end
											endfunction
											for (_gv_block_idx_3 = 0; _gv_block_idx_3 < BLOCK_SIZE; _gv_block_idx_3 = _gv_block_idx_3 + 1) begin : g_blocks
												localparam block_idx = _gv_block_idx_3;
												// Trace: src/VX_dispatch_unit.sv:74:9
												wire [0:0] issue_idx = issue_indices[block_idx+:1];
												// Trace: src/VX_dispatch_unit.sv:75:9
												wire valid_p;
												wire ready_p;
												if (1) begin : g_full_threads
													// Trace: src/VX_dispatch_unit.sv:168:13
													assign valid_p = dispatch_valid[issue_idx];
													// Trace: src/VX_dispatch_unit.sv:169:13
													assign block_tmask[block_idx * 4+:4] = dispatch_data[(issue_idx * 472) + DATA_TMASK_OFF+:4];
													// Trace: src/VX_dispatch_unit.sv:170:13
													assign block_regs[32 * ((block_idx * 3) * 4)+:128] = dispatch_data[(issue_idx * 472) + 256+:128];
													// Trace: src/VX_dispatch_unit.sv:171:13
													assign block_regs[32 * (((block_idx * 3) + 1) * 4)+:128] = dispatch_data[(issue_idx * 472) + 128+:128];
													// Trace: src/VX_dispatch_unit.sv:172:13
													assign block_regs[32 * (((block_idx * 3) + 2) * 4)+:128] = dispatch_data[issue_idx * 472+:128];
													// Trace: src/VX_dispatch_unit.sv:173:13
													assign block_pid[block_idx+:1] = 1'sb0;
													// Trace: src/VX_dispatch_unit.sv:174:13
													assign block_sop[block_idx] = 1'b1;
													// Trace: src/VX_dispatch_unit.sv:175:13
													assign block_eop[block_idx] = 1'b1;
													// Trace: src/VX_dispatch_unit.sv:176:13
													assign block_ready[block_idx] = ready_p;
													// Trace: src/VX_dispatch_unit.sv:177:13
													assign block_done[block_idx] = ready_p || ~valid_p;
												end
												// Trace: src/VX_dispatch_unit.sv:179:9
												wire [0:0] isw;
												if (1) begin : g_isw
													// Trace: src/VX_dispatch_unit.sv:187:13
													assign isw = block_idx;
												end
												// Trace: src/VX_dispatch_unit.sv:189:9
												wire [1:0] block_wid = VX_gpu_pkg_wis_to_wid(dispatch_data[(issue_idx * 472) + 469+:VX_gpu_pkg_ISSUE_WIS_W], isw);
												// Trace: src/VX_dispatch_unit.sv:190:9
												wire [474:0] execute_data;
												reg [474:0] execute_data_w;
												// Trace: src/VX_dispatch_unit.sv:191:9
												VX_elastic_buffer #(
													.DATAW(OUT_DATAW),
													.SIZE(2),
													.OUT_REG(1)
												) buf_out(
													.clk(clk),
													.reset(reset),
													.valid_in(valid_p),
													.ready_in(ready_p),
													.data_in({dispatch_data[(issue_idx * 472) + 471-:1], block_wid, block_tmask[block_idx * 4+:4], dispatch_data[(issue_idx * 472) + 464-:81], block_regs[32 * ((block_idx * 3) * 4)+:128], block_regs[32 * (((block_idx * 3) + 1) * 4)+:128], block_regs[32 * (((block_idx * 3) + 2) * 4)+:128], block_pid[block_idx+:1], block_sop[block_idx], block_eop[block_idx]}),
													.data_out(execute_data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[block_idx + _mbase_execute_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[block_idx + _mbase_execute_if].ready)
												);
												if (1) begin : g_execute_data_w_full
													// Trace: src/VX_dispatch_unit.sv:218:13
													always @(*) begin
														// Trace: src/VX_dispatch_unit.sv:219:17
														execute_data_w = execute_data;
														// Trace: src/VX_dispatch_unit.sv:220:17
														execute_data_w[2:0] = 3'b011;
													end
												end
												// Trace: src/VX_dispatch_unit.sv:223:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[block_idx + _mbase_execute_if].data = execute_data_w;
											end
											// Trace: src/VX_dispatch_unit.sv:225:5
											reg [0:0] ready_in;
											// Trace: src/VX_dispatch_unit.sv:226:5
											always @(*) begin
												// Trace: src/VX_dispatch_unit.sv:227:9
												ready_in = 0;
												// Trace: src/VX_dispatch_unit.sv:228:9
												begin : sv2v_autoblock_18
													// Trace: src/VX_dispatch_unit.sv:228:14
													integer block_idx;
													// Trace: src/VX_dispatch_unit.sv:228:14
													for (block_idx = 0; block_idx < BLOCK_SIZE; block_idx = block_idx + 1)
														begin
															// Trace: src/VX_dispatch_unit.sv:229:13
															ready_in[issue_indices[block_idx+:1]] = block_ready[block_idx] && block_eop[block_idx];
														end
												end
											end
											// Trace: src/VX_dispatch_unit.sv:232:5
											assign dispatch_ready = ready_in;
										end
										assign dispatch_unit.clk = clk;
										assign dispatch_unit.reset = reset;
										// Trace: src/VX_sfu_unit.sv:37:5
										// expanded interface instance: pe_execute_if
										localparam _param_C9035_NUM_LANES = NUM_LANES;
										genvar _arr_C9035;
										for (_arr_C9035 = 0; _arr_C9035 <= 1; _arr_C9035 = _arr_C9035 + 1) begin : pe_execute_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_execute_if.sv:2:15
											localparam NUM_LANES = _param_C9035_NUM_LANES;
											// Trace: src/VX_execute_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_execute_if.sv:5:5
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_execute_if.sv:22:5
											wire valid;
											// Trace: src/VX_execute_if.sv:23:5
											wire [474:0] data;
											// Trace: src/VX_execute_if.sv:24:5
											wire ready;
											// Trace: src/VX_execute_if.sv:25:5
											// Trace: src/VX_execute_if.sv:30:5
										end
										// Trace: src/VX_sfu_unit.sv:40:5
										// expanded interface instance: pe_commit_if
										localparam _param_0FC39_NUM_LANES = NUM_LANES;
										genvar _arr_0FC39;
										for (_arr_0FC39 = 0; _arr_0FC39 <= 1; _arr_0FC39 = _arr_0FC39 + 1) begin : pe_commit_if
											// Trace: src/VX_commit_if.sv:2:15
											localparam NUM_LANES = _param_0FC39_NUM_LANES;
											// Trace: src/VX_commit_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_commit_if.sv:5:5
											// removed localparam type data_t
											// Trace: src/VX_commit_if.sv:17:5
											wire valid;
											// Trace: src/VX_commit_if.sv:18:5
											wire [175:0] data;
											// Trace: src/VX_commit_if.sv:19:5
											wire ready;
											// Trace: src/VX_commit_if.sv:20:5
											// Trace: src/VX_commit_if.sv:25:5
										end
										// Trace: src/VX_sfu_unit.sv:43:5
										reg [0:0] pe_select;
										// Trace: src/VX_sfu_unit.sv:44:5
										always @(*) begin
											// Trace: src/VX_sfu_unit.sv:45:9
											pe_select = PE_IDX_WCTL;
											// Trace: src/VX_sfu_unit.sv:46:9
											if ((per_block_execute_if[0].data[436-:4] >= 6) && (per_block_execute_if[0].data[436-:4] <= 8))
												// Trace: src/VX_sfu_unit.sv:47:13
												pe_select = PE_IDX_CSRS;
										end
										// Trace: src/VX_sfu_unit.sv:49:5
										// expanded module instance: pe_switch
										localparam _bbase_3D12E_execute_in_if = 0;
										localparam _bbase_3D12E_commit_out_if = 0;
										localparam _bbase_3D12E_execute_out_if = 0;
										localparam _bbase_3D12E_commit_in_if = 0;
										localparam _param_3D12E_PE_COUNT = PE_COUNT;
										localparam _param_3D12E_NUM_LANES = NUM_LANES;
										localparam _param_3D12E_ARBITER = "R";
										localparam _param_3D12E_REQ_OUT_BUF = 0;
										localparam _param_3D12E_RSP_OUT_BUF = 3;
										if (1) begin : pe_switch
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_pe_switch.sv:2:15
											localparam PE_COUNT = _param_3D12E_PE_COUNT;
											// Trace: src/VX_pe_switch.sv:3:15
											localparam NUM_LANES = _param_3D12E_NUM_LANES;
											// Trace: src/VX_pe_switch.sv:4:15
											localparam REQ_OUT_BUF = _param_3D12E_REQ_OUT_BUF;
											// Trace: src/VX_pe_switch.sv:5:15
											localparam RSP_OUT_BUF = _param_3D12E_RSP_OUT_BUF;
											// Trace: src/VX_pe_switch.sv:6:16
											localparam ARBITER = _param_3D12E_ARBITER;
											// Trace: src/VX_pe_switch.sv:7:15
											localparam PE_SEL_BITS = 1;
											// Trace: src/VX_pe_switch.sv:9:5
											wire clk;
											// Trace: src/VX_pe_switch.sv:10:5
											wire reset;
											// Trace: src/VX_pe_switch.sv:11:5
											wire [0:0] pe_sel;
											// Trace: src/VX_pe_switch.sv:12:5
											localparam _mbase_execute_in_if = _bbase_3D12E_execute_in_if;
											// Trace: src/VX_pe_switch.sv:13:5
											localparam _mbase_commit_out_if = _bbase_3D12E_commit_out_if;
											// Trace: src/VX_pe_switch.sv:14:5
											localparam _mbase_execute_out_if = 0;
											// Trace: src/VX_pe_switch.sv:15:5
											localparam _mbase_commit_in_if = 0;
											// Trace: src/VX_pe_switch.sv:17:5
											localparam PID_BITS = 0;
											// Trace: src/VX_pe_switch.sv:18:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_pe_switch.sv:19:5
											// removed localparam type VX_gpu_pkg_alu_args_t
											// removed localparam type VX_gpu_pkg_csr_args_t
											// removed localparam type VX_gpu_pkg_fpu_args_t
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											localparam REQ_DATAW = 475;
											// Trace: src/VX_pe_switch.sv:20:5
											localparam RSP_DATAW = 176;
											// Trace: src/VX_pe_switch.sv:21:5
											wire [1:0] pe_req_valid;
											// Trace: src/VX_pe_switch.sv:22:5
											wire [949:0] pe_req_data;
											// Trace: src/VX_pe_switch.sv:23:5
											wire [1:0] pe_req_ready;
											// Trace: src/VX_pe_switch.sv:24:5
											VX_stream_switch #(
												.DATAW(REQ_DATAW),
												.NUM_INPUTS(1),
												.NUM_OUTPUTS(PE_COUNT),
												.OUT_BUF(REQ_OUT_BUF)
											) req_switch(
												.clk(clk),
												.reset(reset),
												.sel_in(pe_sel),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[_mbase_execute_in_if].valid),
												.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[_mbase_execute_in_if].ready),
												.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[_mbase_execute_in_if].data),
												.data_out(pe_req_data),
												.valid_out(pe_req_valid),
												.ready_out(pe_req_ready)
											);
											// Trace: src/VX_pe_switch.sv:40:5
											genvar _gv_i_14;
											for (_gv_i_14 = 0; _gv_i_14 < PE_COUNT; _gv_i_14 = _gv_i_14 + 1) begin : g_execute_out_if
												localparam i = _gv_i_14;
												// Trace: src/VX_pe_switch.sv:41:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[i + _mbase_execute_out_if].valid = pe_req_valid[i];
												// Trace: src/VX_pe_switch.sv:42:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[i + _mbase_execute_out_if].data = pe_req_data[i * 475+:475];
												// Trace: src/VX_pe_switch.sv:43:9
												assign pe_req_ready[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[i + _mbase_execute_out_if].ready;
											end
											// Trace: src/VX_pe_switch.sv:45:5
											wire [1:0] pe_rsp_valid;
											// Trace: src/VX_pe_switch.sv:46:5
											wire [351:0] pe_rsp_data;
											// Trace: src/VX_pe_switch.sv:47:5
											wire [1:0] pe_rsp_ready;
											// Trace: src/VX_pe_switch.sv:48:5
											genvar _gv_i_15;
											for (_gv_i_15 = 0; _gv_i_15 < PE_COUNT; _gv_i_15 = _gv_i_15 + 1) begin : g_commit_in_if
												localparam i = _gv_i_15;
												// Trace: src/VX_pe_switch.sv:49:9
												assign pe_rsp_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[i + _mbase_commit_in_if].valid;
												// Trace: src/VX_pe_switch.sv:50:9
												assign pe_rsp_data[i * 176+:176] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[i + _mbase_commit_in_if].data;
												// Trace: src/VX_pe_switch.sv:51:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[i + _mbase_commit_in_if].ready = pe_rsp_ready[i];
											end
											// Trace: src/VX_pe_switch.sv:53:5
											VX_stream_arb #(
												.NUM_INPUTS(PE_COUNT),
												.DATAW(RSP_DATAW),
												.ARBITER(ARBITER),
												.OUT_BUF(RSP_OUT_BUF)
											) rsp_arb(
												.clk(clk),
												.reset(reset),
												.valid_in(pe_rsp_valid),
												.ready_in(pe_rsp_ready),
												.data_in(pe_rsp_data),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_commit_if[_mbase_commit_out_if].data),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_commit_if[_mbase_commit_out_if].valid),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_commit_if[_mbase_commit_out_if].ready),
												.sel_out()
											);
										end
										assign pe_switch.clk = clk;
										assign pe_switch.reset = reset;
										assign pe_switch.pe_sel = pe_select;
										// Trace: src/VX_sfu_unit.sv:64:5
										// expanded module instance: wctl_unit
										localparam _bbase_F22EA_execute_if = PE_IDX_WCTL;
										localparam _bbase_F22EA_commit_if = PE_IDX_WCTL;
										localparam _param_F22EA_INSTANCE_ID = "";
										localparam _param_F22EA_NUM_LANES = NUM_LANES;
										if (1) begin : wctl_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_wctl_unit.sv:2:16
											localparam INSTANCE_ID = _param_F22EA_INSTANCE_ID;
											// Trace: src/VX_wctl_unit.sv:3:15
											localparam NUM_LANES = _param_F22EA_NUM_LANES;
											// Trace: src/VX_wctl_unit.sv:5:5
											wire clk;
											// Trace: src/VX_wctl_unit.sv:6:5
											wire reset;
											// Trace: src/VX_wctl_unit.sv:7:5
											localparam _mbase_execute_if = _bbase_F22EA_execute_if;
											// Trace: src/VX_wctl_unit.sv:8:5
											// removed modport instance warp_ctl_if
											// Trace: src/VX_wctl_unit.sv:9:5
											localparam _mbase_commit_if = _bbase_F22EA_commit_if;
											// Trace: src/VX_wctl_unit.sv:11:5
											localparam LANE_BITS = 2;
											// Trace: src/VX_wctl_unit.sv:12:5
											localparam PID_BITS = 0;
											// Trace: src/VX_wctl_unit.sv:13:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_wctl_unit.sv:14:5
											// removed localparam type VX_gpu_pkg_barrier_t
											// removed localparam type VX_gpu_pkg_join_t
											// removed localparam type VX_gpu_pkg_split_t
											// removed localparam type VX_gpu_pkg_tmc_t
											// removed localparam type VX_gpu_pkg_wspawn_t
											localparam WCTL_WIDTH = 91;
											// Trace: src/VX_wctl_unit.sv:15:5
											localparam DATAW = 141;
											// Trace: src/VX_wctl_unit.sv:16:5
											wire [4:0] tmc;
											wire [4:0] tmc_r;
											// Trace: src/VX_wctl_unit.sv:17:5
											wire [35:0] wspawn;
											wire [35:0] wspawn_r;
											// Trace: src/VX_wctl_unit.sv:18:5
											wire [40:0] split;
											wire [40:0] split_r;
											// Trace: src/VX_wctl_unit.sv:19:5
											wire [2:0] sjoin;
											wire [2:0] sjoin_r;
											// Trace: src/VX_wctl_unit.sv:20:5
											wire [5:0] barrier;
											wire [5:0] barrier_r;
											// Trace: src/VX_wctl_unit.sv:21:5
											wire is_wspawn = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[436-:4] == 4'h1;
											// Trace: src/VX_wctl_unit.sv:22:5
											wire is_tmc = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[436-:4] == 4'h0;
											// Trace: src/VX_wctl_unit.sv:23:5
											wire is_pred = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[436-:4] == 4'h5;
											// Trace: src/VX_wctl_unit.sv:24:5
											wire is_split = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[436-:4] == 4'h2;
											// Trace: src/VX_wctl_unit.sv:25:5
											wire is_join = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[436-:4] == 4'h3;
											// Trace: src/VX_wctl_unit.sv:26:5
											wire is_bar = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[436-:4] == 4'h4;
											// Trace: src/VX_wctl_unit.sv:27:5
											wire [1:0] tid;
											// Trace: src/VX_wctl_unit.sv:28:5
											if (1) begin : g_tid
												// Trace: src/VX_wctl_unit.sv:29:9
												assign tid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[387+:LANE_BITS];
											end
											// Trace: src/VX_wctl_unit.sv:33:5
											wire [31:0] rs1_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[259 + (tid * 32)+:32];
											// Trace: src/VX_wctl_unit.sv:34:5
											wire [31:0] rs2_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[131 + (tid * 32)+:32];
											// Trace: src/VX_wctl_unit.sv:35:5
											wire not_pred = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[396];
											// Trace: src/VX_wctl_unit.sv:36:5
											wire [3:0] taken;
											// Trace: src/VX_wctl_unit.sv:37:5
											genvar _gv_i_16;
											for (_gv_i_16 = 0; _gv_i_16 < NUM_LANES; _gv_i_16 = _gv_i_16 + 1) begin : g_taken
												localparam i = _gv_i_16;
												// Trace: src/VX_wctl_unit.sv:38:9
												assign taken[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[259 + (i * 32)] ^ not_pred;
											end
											// Trace: src/VX_wctl_unit.sv:40:5
											reg [3:0] then_tmask_r;
											reg [3:0] then_tmask_n;
											// Trace: src/VX_wctl_unit.sv:41:5
											reg [3:0] else_tmask_r;
											reg [3:0] else_tmask_n;
											// Trace: src/VX_wctl_unit.sv:42:5
											always @(*) begin
												// Trace: src/VX_wctl_unit.sv:43:9
												then_tmask_n = then_tmask_r;
												// Trace: src/VX_wctl_unit.sv:44:9
												else_tmask_n = else_tmask_r;
												// Trace: src/VX_wctl_unit.sv:45:9
												if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[1]) begin
													// Trace: src/VX_wctl_unit.sv:46:13
													then_tmask_n = 1'sb0;
													// Trace: src/VX_wctl_unit.sv:47:13
													else_tmask_n = 1'sb0;
												end
												// Trace: src/VX_wctl_unit.sv:49:9
												then_tmask_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[2] * NUM_LANES+:NUM_LANES] = taken & Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[471-:4];
												// Trace: src/VX_wctl_unit.sv:50:9
												else_tmask_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[2] * NUM_LANES+:NUM_LANES] = ~taken & Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[471-:4];
											end
											// Trace: src/VX_wctl_unit.sv:52:5
											always @(posedge clk)
												// Trace: src/VX_wctl_unit.sv:53:9
												if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].valid) begin
													// Trace: src/VX_wctl_unit.sv:54:13
													then_tmask_r <= then_tmask_n;
													// Trace: src/VX_wctl_unit.sv:55:13
													else_tmask_r <= else_tmask_n;
												end
											// Trace: src/VX_wctl_unit.sv:58:5
											wire has_then = then_tmask_n != 0;
											// Trace: src/VX_wctl_unit.sv:59:5
											wire has_else = else_tmask_n != 0;
											// Trace: src/VX_wctl_unit.sv:60:5
											wire [3:0] pred_mask = (has_then ? then_tmask_n : rs2_data[3:0]);
											// Trace: src/VX_wctl_unit.sv:61:5
											assign tmc[4] = is_tmc || is_pred;
											// Trace: src/VX_wctl_unit.sv:62:5
											assign tmc[3-:4] = (is_pred ? pred_mask : rs1_data[3:0]);
											// Trace: src/VX_wctl_unit.sv:63:5
											wire [2:0] then_tmask_cnt;
											wire [2:0] else_tmask_cnt;
											// Trace: src/VX_wctl_unit.sv:64:5
											VX_popcount #(
												.N(4),
												.MODEL(1)
											) __then_tmask_cnt__(
												.data_in(then_tmask_n),
												.data_out(then_tmask_cnt)
											);
											// Trace: src/VX_wctl_unit.sv:71:5
											VX_popcount #(
												.N(4),
												.MODEL(1)
											) __else_tmask_cnt__(
												.data_in(else_tmask_n),
												.data_out(else_tmask_cnt)
											);
											// Trace: src/VX_wctl_unit.sv:78:5
											wire then_first = then_tmask_cnt >= else_tmask_cnt;
											// Trace: src/VX_wctl_unit.sv:79:5
											wire [3:0] taken_tmask = (then_first ? then_tmask_n : else_tmask_n);
											// Trace: src/VX_wctl_unit.sv:80:5
											wire [3:0] ntaken_tmask = (then_first ? else_tmask_n : then_tmask_n);
											// Trace: src/VX_wctl_unit.sv:81:5
											assign split[40] = is_split;
											// Trace: src/VX_wctl_unit.sv:82:5
											assign split[39] = has_then && has_else;
											// Trace: src/VX_wctl_unit.sv:83:5
											assign split[38-:4] = taken_tmask;
											// Trace: src/VX_wctl_unit.sv:84:5
											assign split[34-:4] = ntaken_tmask;
											// Trace: src/VX_wctl_unit.sv:85:5
											assign split[30-:31] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[467-:31] + 31'sd2;
											// Trace: src/VX_wctl_unit.sv:86:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.dvstack_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[473-:2];
											// Trace: src/VX_wctl_unit.sv:87:5
											wire [1:0] dvstack_ptr;
											// Trace: src/VX_wctl_unit.sv:88:5
											assign sjoin[2] = is_join;
											// Trace: src/VX_wctl_unit.sv:89:5
											assign sjoin[1-:2] = rs1_data[1:0];
											// Trace: src/VX_wctl_unit.sv:90:5
											assign barrier[5] = is_bar;
											// Trace: src/VX_wctl_unit.sv:91:5
											assign barrier[4-:1] = rs1_data[0:0];
											// Trace: src/VX_wctl_unit.sv:92:5
											assign barrier[3] = 1'b0;
											// Trace: src/VX_wctl_unit.sv:93:5
											assign barrier[2-:2] = rs2_data[1:0] - sv2v_cast_2C231_signed(1);
											// Trace: src/VX_wctl_unit.sv:94:5
											assign barrier[0] = rs2_data[1:0] == sv2v_cast_2C231_signed(1);
											// Trace: src/VX_wctl_unit.sv:95:5
											wire [3:0] wspawn_wmask;
											// Trace: src/VX_wctl_unit.sv:96:5
											genvar _gv_i_17;
											for (_gv_i_17 = 0; _gv_i_17 < 4; _gv_i_17 = _gv_i_17 + 1) begin : g_wspawn_wmask
												localparam i = _gv_i_17;
												// Trace: src/VX_wctl_unit.sv:97:9
												assign wspawn_wmask[i] = (i < rs1_data[2:0]) && (i != Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[473-:2]);
											end
											// Trace: src/VX_wctl_unit.sv:99:5
											assign wspawn[35] = is_wspawn;
											// Trace: src/VX_wctl_unit.sv:100:5
											assign wspawn[34-:4] = wspawn_wmask;
											// Trace: src/VX_wctl_unit.sv:101:5
											assign wspawn[30-:31] = rs2_data[1+:31];
											// Trace: src/VX_wctl_unit.sv:102:5
											VX_elastic_buffer #(
												.DATAW(DATAW),
												.SIZE(2)
											) rsp_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].valid),
												.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].ready),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[474], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[473-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[471-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[467-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[394-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[395], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[0], tmc, wspawn, split, sjoin, barrier, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.dvstack_ptr}),
												.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[175], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[174-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[172-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[168-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[136-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[137], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[0], tmc_r, wspawn_r, split_r, sjoin_r, barrier_r, dvstack_ptr}),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].valid),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].ready)
											);
											// Trace: src/VX_wctl_unit.sv:115:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].ready) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[0];
											// Trace: src/VX_wctl_unit.sv:116:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[174-:2];
											// Trace: src/VX_wctl_unit.sv:117:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.tmc = tmc_r;
											// Trace: src/VX_wctl_unit.sv:118:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wspawn = wspawn_r;
											// Trace: src/VX_wctl_unit.sv:119:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split = split_r;
											// Trace: src/VX_wctl_unit.sv:120:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.sjoin = sjoin_r;
											// Trace: src/VX_wctl_unit.sv:121:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier = barrier_r;
											// Trace: src/VX_wctl_unit.sv:122:5
											genvar _gv_i_18;
											for (_gv_i_18 = 0; _gv_i_18 < NUM_LANES; _gv_i_18 = _gv_i_18 + 1) begin : g_commit_if
												localparam i = _gv_i_18;
												// Trace: src/VX_wctl_unit.sv:123:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[3 + (i * 32)+:32] = sv2v_cast_32(dvstack_ptr);
											end
										end
										assign wctl_unit.clk = clk;
										assign wctl_unit.reset = reset;
										// Trace: src/VX_sfu_unit.sv:74:5
										// expanded module instance: csr_unit
										localparam _bbase_BED2E_execute_if = PE_IDX_CSRS;
										localparam _bbase_BED2E_fpu_csr_if = 0;
										localparam _bbase_BED2E_commit_if = PE_IDX_CSRS;
										localparam _param_BED2E_INSTANCE_ID = "";
										localparam _param_BED2E_CORE_ID = CORE_ID;
										localparam _param_BED2E_NUM_LANES = NUM_LANES;
										if (1) begin : csr_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_csr_unit.sv:2:16
											localparam INSTANCE_ID = _param_BED2E_INSTANCE_ID;
											// Trace: src/VX_csr_unit.sv:3:15
											localparam CORE_ID = _param_BED2E_CORE_ID;
											// Trace: src/VX_csr_unit.sv:4:15
											localparam NUM_LANES = _param_BED2E_NUM_LANES;
											// Trace: src/VX_csr_unit.sv:6:5
											wire clk;
											// Trace: src/VX_csr_unit.sv:7:5
											wire reset;
											// Trace: src/VX_csr_unit.sv:8:5
											// removed localparam type VX_gpu_pkg_base_dcrs_t
											wire [71:0] base_dcrs;
											// Trace: src/VX_csr_unit.sv:9:5
											localparam _mbase_fpu_csr_if = 0;
											// Trace: src/VX_csr_unit.sv:10:5
											// removed modport instance commit_csr_if
											// Trace: src/VX_csr_unit.sv:11:5
											// removed modport instance sched_csr_if
											// Trace: src/VX_csr_unit.sv:12:5
											localparam _mbase_execute_if = _bbase_BED2E_execute_if;
											// Trace: src/VX_csr_unit.sv:13:5
											localparam _mbase_commit_if = _bbase_BED2E_commit_if;
											// Trace: src/VX_csr_unit.sv:15:5
											localparam PID_BITS = 0;
											// Trace: src/VX_csr_unit.sv:16:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_csr_unit.sv:17:5
											localparam DATAW = 176;
											// Trace: src/VX_csr_unit.sv:18:5
											reg [127:0] csr_read_data;
											// Trace: src/VX_csr_unit.sv:19:5
											reg [31:0] csr_write_data;
											// Trace: src/VX_csr_unit.sv:20:5
											wire [31:0] csr_read_data_ro;
											wire [31:0] csr_read_data_rw;
											// Trace: src/VX_csr_unit.sv:21:5
											wire [31:0] csr_req_data;
											// Trace: src/VX_csr_unit.sv:22:5
											reg csr_rd_enable;
											// Trace: src/VX_csr_unit.sv:23:5
											wire csr_wr_enable;
											// Trace: src/VX_csr_unit.sv:24:5
											wire csr_req_ready;
											// Trace: src/VX_csr_unit.sv:25:5
											wire [11:0] csr_addr = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[412-:12];
											// Trace: src/VX_csr_unit.sv:26:5
											wire [4:0] csr_imm = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[400-:5];
											// Trace: src/VX_csr_unit.sv:27:5
											wire is_fpu_csr = csr_addr <= 12'h003;
											// Trace: src/VX_csr_unit.sv:28:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.alm_empty_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[473-:2];
											// Trace: src/VX_csr_unit.sv:29:5
											wire no_pending_instr = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.alm_empty || ~is_fpu_csr;
											// Trace: src/VX_csr_unit.sv:30:5
											wire csr_req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].valid && no_pending_instr;
											// Trace: src/VX_csr_unit.sv:31:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].ready = csr_req_ready && no_pending_instr;
											// Trace: src/VX_csr_unit.sv:32:5
											wire [127:0] rs1_data;
											// Trace: src/VX_csr_unit.sv:33:5
											genvar _gv_i_191;
											for (_gv_i_191 = 0; _gv_i_191 < NUM_LANES; _gv_i_191 = _gv_i_191 + 1) begin : g_rs1_data
												localparam i = _gv_i_191;
												// Trace: src/VX_csr_unit.sv:34:9
												assign rs1_data[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[259 + (i * 32)+:32];
											end
											// Trace: src/VX_csr_unit.sv:36:5
											wire csr_write_enable = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[436-:4] == 4'h6;
											// Trace: src/VX_csr_unit.sv:37:5
											// expanded module instance: csr_data
											localparam _bbase_9D0B6_fpu_csr_if = 0;
											localparam _param_9D0B6_INSTANCE_ID = INSTANCE_ID;
											localparam _param_9D0B6_CORE_ID = CORE_ID;
											if (1) begin : csr_data
												// removed import VX_gpu_pkg::*;
												// removed import VX_fpu_pkg::*;
												// Trace: src/VX_csr_data.sv:5:16
												localparam INSTANCE_ID = _param_9D0B6_INSTANCE_ID;
												// Trace: src/VX_csr_data.sv:6:15
												localparam CORE_ID = _param_9D0B6_CORE_ID;
												// Trace: src/VX_csr_data.sv:8:5
												wire clk;
												// Trace: src/VX_csr_data.sv:9:5
												wire reset;
												// Trace: src/VX_csr_data.sv:10:5
												// removed localparam type VX_gpu_pkg_base_dcrs_t
												wire [71:0] base_dcrs;
												// Trace: src/VX_csr_data.sv:11:5
												// removed modport instance commit_csr_if
												// Trace: src/VX_csr_data.sv:12:5
												localparam _mbase_fpu_csr_if = 0;
												// Trace: src/VX_csr_data.sv:13:5
												wire [43:0] cycles;
												// Trace: src/VX_csr_data.sv:14:5
												wire [3:0] active_warps;
												// Trace: src/VX_csr_data.sv:15:5
												wire [15:0] thread_masks;
												// Trace: src/VX_csr_data.sv:16:5
												wire read_enable;
												// Trace: src/VX_csr_data.sv:17:5
												wire [0:0] read_uuid;
												// Trace: src/VX_csr_data.sv:18:5
												wire [1:0] read_wid;
												// Trace: src/VX_csr_data.sv:19:5
												wire [11:0] read_addr;
												// Trace: src/VX_csr_data.sv:20:5
												wire [31:0] read_data_ro;
												// Trace: src/VX_csr_data.sv:21:5
												wire [31:0] read_data_rw;
												// Trace: src/VX_csr_data.sv:22:5
												wire write_enable;
												// Trace: src/VX_csr_data.sv:23:5
												wire [0:0] write_uuid;
												// Trace: src/VX_csr_data.sv:24:5
												wire [1:0] write_wid;
												// Trace: src/VX_csr_data.sv:25:5
												wire [11:0] write_addr;
												// Trace: src/VX_csr_data.sv:26:5
												wire [31:0] write_data;
												// Trace: src/VX_csr_data.sv:28:5
												reg [31:0] mscratch;
												// Trace: src/VX_csr_data.sv:29:5
												// removed localparam type VX_fpu_pkg_fflags_t
												reg [31:0] fcsr;
												reg [31:0] fcsr_n;
												// Trace: src/VX_csr_data.sv:30:5
												wire [0:0] fpu_write_enable;
												// Trace: src/VX_csr_data.sv:31:5
												wire [1:0] fpu_write_wid;
												// Trace: src/VX_csr_data.sv:32:5
												wire [4:0] fpu_write_fflags;
												// Trace: src/VX_csr_data.sv:33:5
												genvar _gv_i_44;
												for (_gv_i_44 = 0; _gv_i_44 < 1; _gv_i_44 = _gv_i_44 + 1) begin : g_fpu_write
													localparam i = _gv_i_44;
													// Trace: src/VX_csr_data.sv:34:9
													assign fpu_write_enable[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[i + _mbase_fpu_csr_if].write_enable;
													// Trace: src/VX_csr_data.sv:35:9
													assign fpu_write_wid[i * 2+:2] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[i + _mbase_fpu_csr_if].write_wid;
													// Trace: src/VX_csr_data.sv:36:9
													assign fpu_write_fflags[i * 5+:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[i + _mbase_fpu_csr_if].write_fflags;
												end
												// Trace: src/VX_csr_data.sv:38:5
												always @(*) begin
													// Trace: src/VX_csr_data.sv:39:9
													fcsr_n = fcsr;
													// Trace: src/VX_csr_data.sv:40:9
													begin : sv2v_autoblock_19
														// Trace: src/VX_csr_data.sv:40:14
														integer i;
														// Trace: src/VX_csr_data.sv:40:14
														for (i = 0; i < 1; i = i + 1)
															begin
																// Trace: src/VX_csr_data.sv:41:13
																if (fpu_write_enable[i])
																	// Trace: src/VX_csr_data.sv:42:17
																	fcsr_n[(fpu_write_wid[i * 2+:2] * 8) + 4-:5] = fcsr[(fpu_write_wid[i * 2+:2] * 8) + 4-:5] | fpu_write_fflags[i * 5+:5];
															end
													end
													if (write_enable)
														// Trace: src/VX_csr_data.sv:47:13
														case (write_addr)
															12'h001:
																// Trace: src/VX_csr_data.sv:48:26
																fcsr_n[(write_wid * 8) + 4-:5] = write_data[4:0];
															12'h002:
																// Trace: src/VX_csr_data.sv:49:29
																fcsr_n[(write_wid * 8) + 7-:3] = write_data[2:0];
															12'h003:
																// Trace: src/VX_csr_data.sv:50:28
																fcsr_n[write_wid * 8+:8] = write_data[7:0];
															default:
																;
														endcase
												end
												// Trace: src/VX_csr_data.sv:55:5
												genvar _gv_i_45;
												for (_gv_i_45 = 0; _gv_i_45 < 1; _gv_i_45 = _gv_i_45 + 1) begin : g_fpu_csr_read_frm
													localparam i = _gv_i_45;
													// Trace: src/VX_csr_data.sv:56:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[i + _mbase_fpu_csr_if].read_frm = fcsr[(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.fpu_csr_if[i + _mbase_fpu_csr_if].read_wid * 8) + 7-:3];
												end
												// Trace: src/VX_csr_data.sv:58:5
												always @(posedge clk)
													// Trace: src/VX_csr_data.sv:59:9
													if (reset)
														// Trace: src/VX_csr_data.sv:60:13
														fcsr <= 1'sb0;
													else
														// Trace: src/VX_csr_data.sv:62:13
														fcsr <= fcsr_n;
												// Trace: src/VX_csr_data.sv:65:5
												always @(posedge clk) begin
													// Trace: src/VX_csr_data.sv:66:9
													if (reset)
														// Trace: src/VX_csr_data.sv:67:13
														mscratch <= base_dcrs[39-:32];
													if (write_enable)
														// Trace: src/VX_csr_data.sv:70:13
														case (write_addr)
															12'h001, 12'h002, 12'h003, 12'h180, 12'h300, 12'h744, 12'h302, 12'h303, 12'h304, 12'h305, 12'h341, 12'h3a0, 12'h3b0:
																;
															12'h340:
																// Trace: src/VX_csr_data.sv:86:21
																mscratch <= write_data;
															default:
																;
														endcase
												end
												// Trace: src/VX_csr_data.sv:94:5
												reg [31:0] read_data_ro_w;
												// Trace: src/VX_csr_data.sv:95:5
												reg [31:0] read_data_rw_w;
												// Trace: src/VX_csr_data.sv:96:5
												reg read_addr_valid_w;
												// Trace: src/VX_csr_data.sv:97:5
												always @(*) begin
													// Trace: src/VX_csr_data.sv:98:9
													read_data_ro_w = 1'sb0;
													// Trace: src/VX_csr_data.sv:99:9
													read_data_rw_w = 1'sb0;
													// Trace: src/VX_csr_data.sv:100:9
													read_addr_valid_w = 1;
													// Trace: src/VX_csr_data.sv:101:9
													case (read_addr)
														12'hf11:
															// Trace: src/VX_csr_data.sv:102:24
															read_data_ro_w = 32'sd0;
														12'hf12:
															// Trace: src/VX_csr_data.sv:103:26
															read_data_ro_w = 32'sd0;
														12'hf13:
															// Trace: src/VX_csr_data.sv:104:27
															read_data_ro_w = 32'sd0;
														12'h301:
															// Trace: src/VX_csr_data.sv:105:29
															read_data_ro_w = 32'h40901120;
														12'h001:
															// Trace: src/VX_csr_data.sv:131:27
															read_data_rw_w = sv2v_cast_32(fcsr[(read_wid * 8) + 4-:5]);
														12'h002:
															// Trace: src/VX_csr_data.sv:132:30
															read_data_rw_w = sv2v_cast_32(fcsr[(read_wid * 8) + 7-:3]);
														12'h003:
															// Trace: src/VX_csr_data.sv:133:29
															read_data_rw_w = sv2v_cast_32(fcsr[read_wid * 8+:8]);
														12'h340:
															// Trace: src/VX_csr_data.sv:134:25
															read_data_rw_w = mscratch;
														12'hcc1:
															// Trace: src/VX_csr_data.sv:135:26
															read_data_ro_w = sv2v_cast_32(read_wid);
														12'hcc2:
															// Trace: src/VX_csr_data.sv:136:26
															read_data_ro_w = sv2v_cast_32_signed(CORE_ID);
														12'hcc4:
															// Trace: src/VX_csr_data.sv:137:22
															read_data_ro_w = sv2v_cast_32(thread_masks[read_wid * 4+:4]);
														12'hcc3:
															// Trace: src/VX_csr_data.sv:138:22
															read_data_ro_w = sv2v_cast_32(active_warps);
														12'hfc0:
															// Trace: src/VX_csr_data.sv:139:22
															read_data_ro_w = 32'sd4;
														12'hfc1:
															// Trace: src/VX_csr_data.sv:140:24
															read_data_ro_w = 32'sd4;
														12'hfc2:
															// Trace: src/VX_csr_data.sv:141:24
															read_data_ro_w = 32'sd1;
														12'hfc3:
															// Trace: src/VX_csr_data.sv:142:22
															read_data_ro_w = 32'hffff0000;
														12'hb00:
															// Trace: src/VX_csr_data.sv:143:19
															read_data_ro_w = cycles[31:0];
														12'hb00 + 12'h080:
															// Trace: src/VX_csr_data.sv:144:26
															read_data_ro_w = sv2v_cast_32(cycles[43:32]);
														12'hb01:
															// Trace: src/VX_csr_data.sv:145:23
															read_data_ro_w = 1'sbx;
														12'hb81:
															// Trace: src/VX_csr_data.sv:146:23
															read_data_ro_w = 1'sbx;
														12'hb02:
															// Trace: src/VX_csr_data.sv:147:19
															read_data_ro_w = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_csr_if.instret[31:0];
														12'hb02 + 12'h080:
															// Trace: src/VX_csr_data.sv:148:26
															read_data_ro_w = sv2v_cast_32(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_csr_if.instret[43:32]);
														12'h180, 12'h300, 12'h744, 12'h302, 12'h303, 12'h304, 12'h305, 12'h341, 12'h3a0, 12'h3b0:
															// Trace: src/VX_csr_data.sv:158:23
															read_data_ro_w = 32'sd0;
														default: begin
															// Trace: src/VX_csr_data.sv:160:17
															read_addr_valid_w = 0;
															// Trace: src/VX_csr_data.sv:161:17
															if (((read_addr >= 12'hb03) && (read_addr < 2851)) || ((read_addr >= 12'hb83) && (read_addr < 2979)))
																// Trace: src/VX_csr_data.sv:163:21
																read_addr_valid_w = 1;
														end
													endcase
												end
												// Trace: src/VX_csr_data.sv:168:5
												assign read_data_ro = read_data_ro_w;
												// Trace: src/VX_csr_data.sv:169:5
												assign read_data_rw = read_data_rw_w;
											end
											assign csr_data.clk = clk;
											assign csr_data.reset = reset;
											assign csr_data.base_dcrs = base_dcrs;
											assign csr_data.cycles = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.cycles;
											assign csr_data.active_warps = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.active_warps;
											assign csr_data.thread_masks = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.thread_masks;
											assign csr_data.read_enable = csr_req_valid && csr_rd_enable;
											assign csr_data.read_uuid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[474];
											assign csr_data.read_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[473-:2];
											assign csr_data.read_addr = csr_addr;
											assign csr_read_data_ro = csr_data.read_data_ro;
											assign csr_read_data_rw = csr_data.read_data_rw;
											assign csr_data.write_enable = csr_req_valid && csr_wr_enable;
											assign csr_data.write_uuid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[474];
											assign csr_data.write_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[473-:2];
											assign csr_data.write_addr = csr_addr;
											assign csr_data.write_data = csr_write_data;
											// Trace: src/VX_csr_unit.sv:61:5
											wire [127:0] wtid;
											wire [127:0] gtid;
											// Trace: src/VX_csr_unit.sv:62:5
											genvar _gv_i_192;
											for (_gv_i_192 = 0; _gv_i_192 < NUM_LANES; _gv_i_192 = _gv_i_192 + 1) begin : g_wtid
												localparam i = _gv_i_192;
												if (1) begin : g_no_pid
													// Trace: src/VX_csr_unit.sv:66:13
													assign wtid[i * 32+:32] = i;
												end
											end
											// Trace: src/VX_csr_unit.sv:69:5
											genvar _gv_i_193;
											for (_gv_i_193 = 0; _gv_i_193 < NUM_LANES; _gv_i_193 = _gv_i_193 + 1) begin : g_gtid
												localparam i = _gv_i_193;
												// Trace: src/VX_csr_unit.sv:70:9
												assign gtid[i * 32+:32] = ((sv2v_cast_32_signed(CORE_ID) << 4) + (sv2v_cast_32(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[473-:2]) << 2)) + wtid[i * 32+:32];
											end
											// Trace: src/VX_csr_unit.sv:72:5
											always @(*) begin
												// Trace: src/VX_csr_unit.sv:73:9
												csr_rd_enable = 0;
												// Trace: src/VX_csr_unit.sv:74:9
												case (csr_addr)
													12'hcc0:
														// Trace: src/VX_csr_unit.sv:75:19
														csr_read_data = wtid;
													12'hf14:
														// Trace: src/VX_csr_unit.sv:76:21
														csr_read_data = gtid;
													default: begin
														// Trace: src/VX_csr_unit.sv:78:13
														csr_read_data = {NUM_LANES {csr_read_data_ro | csr_read_data_rw}};
														// Trace: src/VX_csr_unit.sv:79:13
														csr_rd_enable = 1;
													end
												endcase
											end
											// Trace: src/VX_csr_unit.sv:83:5
											assign csr_req_data = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[413] ? sv2v_cast_32(csr_imm) : rs1_data[0+:32]);
											// Trace: src/VX_csr_unit.sv:84:5
											assign csr_wr_enable = csr_write_enable || |csr_req_data;
											// Trace: src/VX_csr_unit.sv:85:5
											always @(*)
												// Trace: src/VX_csr_unit.sv:86:9
												case (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[436-:4])
													4'h6:
														// Trace: src/VX_csr_unit.sv:88:17
														csr_write_data = csr_req_data;
													4'h7:
														// Trace: src/VX_csr_unit.sv:91:17
														csr_write_data = csr_read_data_rw | csr_req_data;
													default:
														// Trace: src/VX_csr_unit.sv:94:17
														csr_write_data = csr_read_data_rw & ~csr_req_data;
												endcase
											// Trace: src/VX_csr_unit.sv:98:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.unlock_warp = ((csr_req_valid && csr_req_ready) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[0]) && is_fpu_csr;
											// Trace: src/VX_csr_unit.sv:99:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.unlock_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[473-:2];
											// Trace: src/VX_csr_unit.sv:100:5
											VX_elastic_buffer #(
												.DATAW(DATAW),
												.SIZE(2)
											) rsp_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(csr_req_valid),
												.ready_in(csr_req_ready),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[474], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[473-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[471-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[467-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[394-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[395], csr_read_data, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[0]}),
												.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[175], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[174-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[172-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[168-:31], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[136-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[137], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[130-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].data[0]}),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].valid),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_commit_if[_mbase_commit_if].ready)
											);
										end
										assign csr_unit.clk = clk;
										assign csr_unit.reset = reset;
										assign csr_unit.base_dcrs = base_dcrs;
										// Trace: src/VX_sfu_unit.sv:88:5
										// expanded module instance: gather_unit
										localparam _bbase_8E516_commit_in_if = 0;
										localparam _bbase_8E516_commit_out_if = 2;
										localparam _param_8E516_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_8E516_NUM_LANES = NUM_LANES;
										localparam _param_8E516_OUT_BUF = 3;
										if (1) begin : gather_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_gather_unit.sv:2:15
											localparam BLOCK_SIZE = _param_8E516_BLOCK_SIZE;
											// Trace: src/VX_gather_unit.sv:3:15
											localparam NUM_LANES = _param_8E516_NUM_LANES;
											// Trace: src/VX_gather_unit.sv:4:15
											localparam OUT_BUF = _param_8E516_OUT_BUF;
											// Trace: src/VX_gather_unit.sv:6:5
											wire clk;
											// Trace: src/VX_gather_unit.sv:7:5
											wire reset;
											// Trace: src/VX_gather_unit.sv:8:5
											localparam _mbase_commit_in_if = 0;
											// Trace: src/VX_gather_unit.sv:9:5
											localparam _mbase_commit_out_if = 2;
											// Trace: src/VX_gather_unit.sv:11:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_gather_unit.sv:12:5
											localparam PID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:13:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:14:5
											localparam DATAW = 176;
											// Trace: src/VX_gather_unit.sv:15:5
											localparam DATA_WIS_OFF = 173;
											// Trace: src/VX_gather_unit.sv:16:5
											wire [0:0] commit_in_valid;
											// Trace: src/VX_gather_unit.sv:17:5
											wire [175:0] commit_in_data;
											// Trace: src/VX_gather_unit.sv:18:5
											wire [0:0] commit_in_ready;
											// Trace: src/VX_gather_unit.sv:19:5
											localparam VX_gpu_pkg_ISSUE_ISW = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											wire [0:0] commit_in_isw;
											// Trace: src/VX_gather_unit.sv:20:5
											genvar _gv_i_208;
											for (_gv_i_208 = 0; _gv_i_208 < BLOCK_SIZE; _gv_i_208 = _gv_i_208 + 1) begin : g_commit_in
												localparam i = _gv_i_208;
												// Trace: src/VX_gather_unit.sv:21:9
												assign commit_in_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_commit_if[i + _mbase_commit_in_if].valid;
												// Trace: src/VX_gather_unit.sv:22:9
												assign commit_in_data[i * 176+:176] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_commit_if[i + _mbase_commit_in_if].data;
												// Trace: src/VX_gather_unit.sv:23:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_commit_if[i + _mbase_commit_in_if].ready = commit_in_ready[i];
												if (1) begin : g_commit_in_isw_full
													// Trace: src/VX_gather_unit.sv:31:13
													assign commit_in_isw[i+:1] = sv2v_cast_1_signed(i);
												end
											end
											// Trace: src/VX_gather_unit.sv:34:5
											reg [0:0] commit_out_valid;
											// Trace: src/VX_gather_unit.sv:35:5
											reg [175:0] commit_out_data;
											// Trace: src/VX_gather_unit.sv:36:5
											wire [0:0] commit_out_ready;
											// Trace: src/VX_gather_unit.sv:37:5
											always @(*) begin
												// Trace: src/VX_gather_unit.sv:38:9
												commit_out_valid = 1'sb0;
												// Trace: src/VX_gather_unit.sv:39:9
												begin : sv2v_autoblock_20
													// Trace: src/VX_gather_unit.sv:39:14
													integer i;
													// Trace: src/VX_gather_unit.sv:39:14
													for (i = 0; i < 1; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:40:13
															commit_out_data[i * 176+:176] = 1'sbx;
														end
												end
												begin : sv2v_autoblock_21
													// Trace: src/VX_gather_unit.sv:42:14
													integer i;
													// Trace: src/VX_gather_unit.sv:42:14
													for (i = 0; i < BLOCK_SIZE; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:43:13
															commit_out_valid[commit_in_isw[i+:1]] = commit_in_valid[i];
															// Trace: src/VX_gather_unit.sv:44:13
															commit_out_data[commit_in_isw[i+:1] * 176+:176] = commit_in_data[i * 176+:176];
														end
												end
											end
											// Trace: src/VX_gather_unit.sv:47:5
											genvar _gv_i_209;
											for (_gv_i_209 = 0; _gv_i_209 < BLOCK_SIZE; _gv_i_209 = _gv_i_209 + 1) begin : g_commit_in_ready
												localparam i = _gv_i_209;
												// Trace: src/VX_gather_unit.sv:48:9
												assign commit_in_ready[i] = commit_out_ready[commit_in_isw[i+:1]];
											end
											// Trace: src/VX_gather_unit.sv:50:5
											genvar _gv_i_210;
											for (_gv_i_210 = 0; _gv_i_210 < 1; _gv_i_210 = _gv_i_210 + 1) begin : g_out_bufs
												localparam i = _gv_i_210;
												// Trace: src/VX_gather_unit.sv:51:9
												// expanded interface instance: commit_tmp_if
												localparam _param_C9958_NUM_LANES = NUM_LANES;
												if (1) begin : commit_tmp_if
													// Trace: src/VX_commit_if.sv:2:15
													localparam NUM_LANES = _param_C9958_NUM_LANES;
													// Trace: src/VX_commit_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_commit_if.sv:5:5
													// removed localparam type data_t
													// Trace: src/VX_commit_if.sv:17:5
													wire valid;
													// Trace: src/VX_commit_if.sv:18:5
													wire [175:0] data;
													// Trace: src/VX_commit_if.sv:19:5
													wire ready;
													// Trace: src/VX_commit_if.sv:20:5
													// Trace: src/VX_commit_if.sv:25:5
												end
												// Trace: src/VX_gather_unit.sv:54:9
												VX_elastic_buffer #(
													.DATAW(DATAW),
													.SIZE(2),
													.OUT_REG(1)
												) out_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(commit_out_valid[i]),
													.ready_in(commit_out_ready[i]),
													.data_in(commit_out_data[i * 176+:176]),
													.data_out(commit_tmp_if.data),
													.valid_out(commit_tmp_if.valid),
													.ready_out(commit_tmp_if.ready)
												);
												// Trace: src/VX_gather_unit.sv:68:9
												wire [3:0] commit_tmask_w;
												// Trace: src/VX_gather_unit.sv:69:9
												wire [127:0] commit_data_w;
												if (1) begin : g_commit_data_no_pid
													// Trace: src/VX_gather_unit.sv:80:13
													assign commit_tmask_w = commit_tmp_if.data[172-:4];
													// Trace: src/VX_gather_unit.sv:81:13
													assign commit_data_w = commit_tmp_if.data[130-:128];
												end
												// Trace: src/VX_gather_unit.sv:83:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].valid = commit_tmp_if.valid;
												// Trace: src/VX_gather_unit.sv:84:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].data = {commit_tmp_if.data[175], commit_tmp_if.data[174-:2], commit_tmask_w, commit_tmp_if.data[168-:31], commit_tmp_if.data[137], commit_tmp_if.data[136-:6], commit_data_w, 1'b0, commit_tmp_if.data[1], commit_tmp_if.data[0]};
												// Trace: src/VX_gather_unit.sv:96:9
												assign commit_tmp_if.ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_out_if].ready;
											end
										end
										assign gather_unit.clk = clk;
										assign gather_unit.reset = reset;
									end
									assign sfu_unit.clk = clk;
									assign sfu_unit.reset = reset;
									assign sfu_unit.base_dcrs = base_dcrs;
								end
								assign execute.clk = clk;
								assign execute.reset = reset;
								assign execute.base_dcrs = base_dcrs;
								// Trace: src/VX_core.sv:94:5
								// expanded module instance: commit
								localparam _bbase_D837E_commit_if = 0;
								localparam _bbase_D837E_writeback_if = 0;
								localparam _param_D837E_INSTANCE_ID = "";
								if (1) begin : commit
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_commit.sv:2:16
									localparam INSTANCE_ID = _param_D837E_INSTANCE_ID;
									// Trace: src/VX_commit.sv:4:5
									wire clk;
									// Trace: src/VX_commit.sv:5:5
									wire reset;
									// Trace: src/VX_commit.sv:6:5
									localparam _mbase_commit_if = 0;
									// Trace: src/VX_commit.sv:7:5
									localparam _mbase_writeback_if = 0;
									// Trace: src/VX_commit.sv:8:5
									// removed modport instance commit_csr_if
									// Trace: src/VX_commit.sv:9:5
									// removed modport instance commit_sched_if
									// Trace: src/VX_commit.sv:11:5
									localparam DATAW = 176;
									// Trace: src/VX_commit.sv:12:5
									localparam COMMIT_SIZEW = 3;
									// Trace: src/VX_commit.sv:13:5
									localparam COMMIT_ALL_SIZEW = 3;
									// Trace: src/VX_commit.sv:14:5
									// expanded interface instance: commit_arb_if
									genvar _arr_25972;
									for (_arr_25972 = 0; _arr_25972 <= 0; _arr_25972 = _arr_25972 + 1) begin : commit_arb_if
										// Trace: src/VX_commit_if.sv:2:15
										localparam NUM_LANES = 4;
										// Trace: src/VX_commit_if.sv:3:15
										localparam PID_WIDTH = 1;
										// Trace: src/VX_commit_if.sv:5:5
										// removed localparam type data_t
										// Trace: src/VX_commit_if.sv:17:5
										wire valid;
										// Trace: src/VX_commit_if.sv:18:5
										wire [175:0] data;
										// Trace: src/VX_commit_if.sv:19:5
										wire ready;
										// Trace: src/VX_commit_if.sv:20:5
										// Trace: src/VX_commit_if.sv:25:5
									end
									// Trace: src/VX_commit.sv:15:5
									wire [0:0] per_issue_commit_fire;
									// Trace: src/VX_commit.sv:16:5
									wire [1:0] per_issue_commit_wid;
									// Trace: src/VX_commit.sv:17:5
									wire [3:0] per_issue_commit_tmask;
									// Trace: src/VX_commit.sv:18:5
									wire [0:0] per_issue_commit_eop;
									// Trace: src/VX_commit.sv:19:5
									genvar _gv_i_46;
									for (_gv_i_46 = 0; _gv_i_46 < 1; _gv_i_46 = _gv_i_46 + 1) begin : g_commit_arbs
										localparam i = _gv_i_46;
										// Trace: src/VX_commit.sv:20:9
										wire [3:0] valid_in;
										// Trace: src/VX_commit.sv:21:9
										wire [703:0] data_in;
										// Trace: src/VX_commit.sv:22:9
										wire [3:0] ready_in;
										genvar _gv_j_4;
										for (_gv_j_4 = 0; _gv_j_4 < 4; _gv_j_4 = _gv_j_4 + 1) begin : g_data_in
											localparam j = _gv_j_4;
											// Trace: src/VX_commit.sv:24:13
											assign valid_in[j] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[((j * 1) + i) + _mbase_commit_if].valid;
											// Trace: src/VX_commit.sv:25:13
											assign data_in[j * 176+:176] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[((j * 1) + i) + _mbase_commit_if].data;
											// Trace: src/VX_commit.sv:26:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[((j * 1) + i) + _mbase_commit_if].ready = ready_in[j];
										end
										// Trace: src/VX_commit.sv:28:9
										VX_stream_arb #(
											.NUM_INPUTS(4),
											.DATAW(DATAW),
											.ARBITER("P"),
											.OUT_BUF(1)
										) commit_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(valid_in),
											.ready_in(ready_in),
											.data_in(data_in),
											.data_out(commit_arb_if[i].data),
											.valid_out(commit_arb_if[i].valid),
											.ready_out(commit_arb_if[i].ready),
											.sel_out()
										);
										// Trace: src/VX_commit.sv:44:9
										assign per_issue_commit_fire[i] = commit_arb_if[i].valid && commit_arb_if[i].ready;
										// Trace: src/VX_commit.sv:45:9
										assign per_issue_commit_tmask[i * 4+:4] = {4 {per_issue_commit_fire[i]}} & commit_arb_if[i].data[172-:4];
										// Trace: src/VX_commit.sv:46:9
										assign per_issue_commit_wid[i * 2+:2] = commit_arb_if[i].data[174-:2];
										// Trace: src/VX_commit.sv:47:9
										assign per_issue_commit_eop[i] = commit_arb_if[i].data[0];
									end
									// Trace: src/VX_commit.sv:49:5
									wire [2:0] commit_size;
									wire [2:0] commit_size_r;
									// Trace: src/VX_commit.sv:50:5
									wire [2:0] commit_size_all_r;
									wire [2:0] commit_size_all_rr;
									// Trace: src/VX_commit.sv:51:5
									wire commit_fire_any;
									wire commit_fire_any_r;
									wire commit_fire_any_rr;
									// Trace: src/VX_commit.sv:52:5
									assign commit_fire_any = |per_issue_commit_fire;
									// Trace: src/VX_commit.sv:53:5
									genvar _gv_i_47;
									for (_gv_i_47 = 0; _gv_i_47 < 1; _gv_i_47 = _gv_i_47 + 1) begin : g_commit_size
										localparam i = _gv_i_47;
										// Trace: src/VX_commit.sv:54:9
										wire [2:0] count;
										// Trace: src/VX_commit.sv:55:5
										VX_popcount #(
											.N(4),
											.MODEL(1)
										) __count__(
											.data_in(per_issue_commit_tmask[i * 4+:4]),
											.data_out(count)
										);
										// Trace: src/VX_commit.sv:62:9
										assign commit_size[i * 3+:3] = count;
									end
									// Trace: src/VX_commit.sv:64:5
									VX_pipe_register #(
										.DATAW(4),
										.RESETW(1)
									) commit_size_reg1(
										.clk(clk),
										.reset(reset),
										.enable(1'b1),
										.data_in({commit_fire_any, commit_size}),
										.data_out({commit_fire_any_r, commit_size_r})
									);
									// Trace: src/VX_commit.sv:74:5
									VX_reduce #(
										.DATAW_IN(COMMIT_SIZEW),
										.DATAW_OUT(COMMIT_ALL_SIZEW),
										.N(1),
										.OP("+")
									) commit_size_reduce(
										.data_in(commit_size_r),
										.data_out(commit_size_all_r)
									);
									// Trace: src/VX_commit.sv:83:5
									VX_pipe_register #(
										.DATAW(4),
										.RESETW(1)
									) commit_size_reg2(
										.clk(clk),
										.reset(reset),
										.enable(1'b1),
										.data_in({commit_fire_any_r, commit_size_all_r}),
										.data_out({commit_fire_any_rr, commit_size_all_rr})
									);
									// Trace: src/VX_commit.sv:93:5
									reg [43:0] instret;
									// Trace: src/VX_commit.sv:94:5
									always @(posedge clk)
										// Trace: src/VX_commit.sv:95:8
										if (reset)
											// Trace: src/VX_commit.sv:96:13
											instret <= 1'sb0;
										else
											// Trace: src/VX_commit.sv:98:13
											if (commit_fire_any_rr)
												// Trace: src/VX_commit.sv:99:17
												instret <= instret + sv2v_cast_44(commit_size_all_rr);
									// Trace: src/VX_commit.sv:103:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_csr_if.instret = instret;
									// Trace: src/VX_commit.sv:104:5
									reg [3:0] committed_warps;
									// Trace: src/VX_commit.sv:105:5
									always @(*) begin
										// Trace: src/VX_commit.sv:106:9
										committed_warps = 0;
										// Trace: src/VX_commit.sv:107:9
										begin : sv2v_autoblock_22
											// Trace: src/VX_commit.sv:107:14
											integer i;
											// Trace: src/VX_commit.sv:107:14
											for (i = 0; i < 1; i = i + 1)
												begin
													// Trace: src/VX_commit.sv:108:13
													if (per_issue_commit_fire[i] && per_issue_commit_eop[i])
														// Trace: src/VX_commit.sv:109:17
														committed_warps[per_issue_commit_wid[i * 2+:2]] = 1;
												end
										end
									end
									// Trace: src/VX_commit.sv:113:5
									VX_pipe_register #(
										.DATAW(4),
										.RESETW(4)
									) committed_pipe_reg(
										.clk(clk),
										.reset(reset),
										.enable(1'b1),
										.data_in(committed_warps),
										.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_sched_if.committed_warps})
									);
									// Trace: src/VX_commit.sv:123:5
									genvar _gv_i_48;
									localparam VX_gpu_pkg_ISSUE_ISW = 0;
									localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
									localparam VX_gpu_pkg_ISSUE_WIS = 2;
									localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS;
									function [1:0] VX_gpu_pkg_wid_to_wis;
										// Trace: src/VX_gpu_pkg.sv:172:9
										input reg [1:0] wid;
										// Trace: src/VX_gpu_pkg.sv:174:9
										begin
											// Trace: src/VX_gpu_pkg.sv:175:13
											VX_gpu_pkg_wid_to_wis = wid >> VX_gpu_pkg_ISSUE_ISW;
										end
									endfunction
									for (_gv_i_48 = 0; _gv_i_48 < 1; _gv_i_48 = _gv_i_48 + 1) begin : g_writeback
										localparam i = _gv_i_48;
										// Trace: src/VX_commit.sv:124:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].valid = commit_arb_if[i].valid && commit_arb_if[i].data[137];
										// Trace: src/VX_commit.sv:125:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[173] = commit_arb_if[i].data[175];
										// Trace: src/VX_commit.sv:126:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[172-:2] = VX_gpu_pkg_wid_to_wis(commit_arb_if[i].data[174-:2]);
										// Trace: src/VX_commit.sv:127:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[166-:31] = commit_arb_if[i].data[168-:31];
										// Trace: src/VX_commit.sv:128:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[170-:4] = commit_arb_if[i].data[172-:4];
										// Trace: src/VX_commit.sv:129:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[135-:6] = commit_arb_if[i].data[136-:6];
										// Trace: src/VX_commit.sv:130:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[129-:128] = commit_arb_if[i].data[130-:128];
										// Trace: src/VX_commit.sv:131:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[1] = commit_arb_if[i].data[1];
										// Trace: src/VX_commit.sv:132:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[0] = commit_arb_if[i].data[0];
										// Trace: src/VX_commit.sv:133:9
										assign commit_arb_if[i].ready = 1'b1;
									end
								end
								assign commit.clk = clk;
								assign commit.reset = reset;
								// Trace: src/VX_core.sv:104:5
								// expanded module instance: mem_unit
								localparam _bbase_A06D0_lsu_mem_if = 0;
								localparam _bbase_A06D0_dcache_bus_if = core_id * VX_gpu_pkg_DCACHE_NUM_REQS;
								localparam _param_A06D0_INSTANCE_ID = INSTANCE_ID;
								if (1) begin : mem_unit
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_unit.sv:2:16
									localparam INSTANCE_ID = _param_A06D0_INSTANCE_ID;
									// Trace: src/VX_mem_unit.sv:4:5
									wire clk;
									// Trace: src/VX_mem_unit.sv:5:5
									wire reset;
									// Trace: src/VX_mem_unit.sv:6:5
									localparam _mbase_lsu_mem_if = 0;
									// Trace: src/VX_mem_unit.sv:7:5
									localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
									localparam VX_gpu_pkg_LSU_WORD_SIZE = 4;
									localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
									localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
									localparam _mbase_dcache_bus_if = _bbase_A06D0_dcache_bus_if;
									// Trace: src/VX_mem_unit.sv:9:5
									localparam VX_gpu_pkg_LSU_MEM_BATCHES = 1;
									localparam VX_gpu_pkg_LSU_TAG_ID_BITS = 1;
									localparam VX_gpu_pkg_LSU_TAG_WIDTH = 2;
									// expanded interface instance: lsu_dcache_if
									localparam _param_9E566_NUM_LANES = 4;
									localparam _param_9E566_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_9E566_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
									genvar _arr_9E566;
									for (_arr_9E566 = 0; _arr_9E566 <= 0; _arr_9E566 = _arr_9E566 + 1) begin : lsu_dcache_if
										// Trace: src/VX_lsu_mem_if.sv:2:15
										localparam NUM_LANES = _param_9E566_NUM_LANES;
										// Trace: src/VX_lsu_mem_if.sv:3:15
										localparam DATA_SIZE = _param_9E566_DATA_SIZE;
										// Trace: src/VX_lsu_mem_if.sv:4:15
										localparam TAG_WIDTH = _param_9E566_TAG_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:5:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_lsu_mem_if.sv:6:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_lsu_mem_if.sv:7:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_lsu_mem_if.sv:8:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_lsu_mem_if.sv:10:5
										// removed localparam type tag_t
										// Trace: src/VX_lsu_mem_if.sv:14:5
										// removed localparam type req_data_t
										// Trace: src/VX_lsu_mem_if.sv:23:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_lsu_mem_if.sv:28:5
										wire req_valid;
										// Trace: src/VX_lsu_mem_if.sv:29:5
										wire [282:0] req_data;
										// Trace: src/VX_lsu_mem_if.sv:30:5
										wire req_ready;
										// Trace: src/VX_lsu_mem_if.sv:31:5
										wire rsp_valid;
										// Trace: src/VX_lsu_mem_if.sv:32:5
										wire [133:0] rsp_data;
										// Trace: src/VX_lsu_mem_if.sv:33:5
										wire rsp_ready;
										// Trace: src/VX_lsu_mem_if.sv:34:5
										// Trace: src/VX_lsu_mem_if.sv:42:5
									end
									// Trace: src/VX_mem_unit.sv:14:5
									localparam LMEM_ADDR_WIDTH = 12;
									// Trace: src/VX_mem_unit.sv:15:6
									// expanded interface instance: lsu_lmem_if
									localparam _param_B7A65_NUM_LANES = 4;
									localparam _param_B7A65_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_B7A65_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
									genvar _arr_B7A65;
									for (_arr_B7A65 = 0; _arr_B7A65 <= 0; _arr_B7A65 = _arr_B7A65 + 1) begin : lsu_lmem_if
										// Trace: src/VX_lsu_mem_if.sv:2:15
										localparam NUM_LANES = _param_B7A65_NUM_LANES;
										// Trace: src/VX_lsu_mem_if.sv:3:15
										localparam DATA_SIZE = _param_B7A65_DATA_SIZE;
										// Trace: src/VX_lsu_mem_if.sv:4:15
										localparam TAG_WIDTH = _param_B7A65_TAG_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:5:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_lsu_mem_if.sv:6:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_lsu_mem_if.sv:7:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_lsu_mem_if.sv:8:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_lsu_mem_if.sv:10:5
										// removed localparam type tag_t
										// Trace: src/VX_lsu_mem_if.sv:14:5
										// removed localparam type req_data_t
										// Trace: src/VX_lsu_mem_if.sv:23:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_lsu_mem_if.sv:28:5
										wire req_valid;
										// Trace: src/VX_lsu_mem_if.sv:29:5
										wire [282:0] req_data;
										// Trace: src/VX_lsu_mem_if.sv:30:5
										wire req_ready;
										// Trace: src/VX_lsu_mem_if.sv:31:5
										wire rsp_valid;
										// Trace: src/VX_lsu_mem_if.sv:32:5
										wire [133:0] rsp_data;
										// Trace: src/VX_lsu_mem_if.sv:33:5
										wire rsp_ready;
										// Trace: src/VX_lsu_mem_if.sv:34:5
										// Trace: src/VX_lsu_mem_if.sv:42:5
									end
									// Trace: src/VX_mem_unit.sv:20:5
									genvar _gv_i_203;
									for (_gv_i_203 = 0; _gv_i_203 < 1; _gv_i_203 = _gv_i_203 + 1) begin : g_lmem_switches
										localparam i = _gv_i_203;
										// Trace: src/VX_mem_unit.sv:21:9
										// expanded module instance: lmem_switch
										localparam _bbase_5CF86_lsu_in_if = i + _mbase_lsu_mem_if;
										localparam _bbase_5CF86_global_out_if = i;
										localparam _bbase_5CF86_local_out_if = i;
										localparam _param_5CF86_REQ0_OUT_BUF = 1;
										localparam _param_5CF86_REQ1_OUT_BUF = 0;
										localparam _param_5CF86_RSP_OUT_BUF = 1;
										localparam _param_5CF86_ARBITER = "P";
										if (1) begin : lmem_switch
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_lmem_switch.sv:2:15
											localparam REQ0_OUT_BUF = _param_5CF86_REQ0_OUT_BUF;
											// Trace: src/VX_lmem_switch.sv:3:15
											localparam REQ1_OUT_BUF = _param_5CF86_REQ1_OUT_BUF;
											// Trace: src/VX_lmem_switch.sv:4:15
											localparam RSP_OUT_BUF = _param_5CF86_RSP_OUT_BUF;
											// Trace: src/VX_lmem_switch.sv:5:16
											localparam ARBITER = _param_5CF86_ARBITER;
											// Trace: src/VX_lmem_switch.sv:7:5
											wire clk;
											// Trace: src/VX_lmem_switch.sv:8:5
											wire reset;
											// Trace: src/VX_lmem_switch.sv:9:5
											localparam _mbase_lsu_in_if = _bbase_5CF86_lsu_in_if;
											// Trace: src/VX_lmem_switch.sv:10:5
											localparam _mbase_global_out_if = _bbase_5CF86_global_out_if;
											// Trace: src/VX_lmem_switch.sv:11:5
											localparam _mbase_local_out_if = _bbase_5CF86_local_out_if;
											// Trace: src/VX_lmem_switch.sv:13:5
											localparam VX_gpu_pkg_LSU_WORD_SIZE = 4;
											localparam VX_gpu_pkg_LSU_ADDR_WIDTH = 30;
											localparam VX_gpu_pkg_LSU_MEM_BATCHES = 1;
											localparam VX_gpu_pkg_LSU_TAG_ID_BITS = 1;
											localparam VX_gpu_pkg_LSU_TAG_WIDTH = 2;
											localparam REQ_DATAW = 283;
											// Trace: src/VX_lmem_switch.sv:14:5
											localparam RSP_DATAW = 134;
											// Trace: src/VX_lmem_switch.sv:15:5
											wire [3:0] is_addr_local_mask;
											// Trace: src/VX_lmem_switch.sv:16:5
											wire req_global_ready;
											// Trace: src/VX_lmem_switch.sv:17:5
											wire req_local_ready;
											// Trace: src/VX_lmem_switch.sv:18:5
											genvar _gv_i_95;
											for (_gv_i_95 = 0; _gv_i_95 < 4; _gv_i_95 = _gv_i_95 + 1) begin : g_is_addr_local_mask
												localparam i = _gv_i_95;
												// Trace: src/VX_lmem_switch.sv:19:9
												assign is_addr_local_mask[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[2 + ((i * 3) + 2)];
											end
											// Trace: src/VX_lmem_switch.sv:21:5
											wire is_addr_global = |(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[282-:4] & ~is_addr_local_mask);
											// Trace: src/VX_lmem_switch.sv:22:5
											wire is_addr_local = |(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[282-:4] & is_addr_local_mask);
											// Trace: src/VX_lmem_switch.sv:23:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_ready = (req_global_ready && is_addr_global) || (req_local_ready && is_addr_local);
											// Trace: src/VX_lmem_switch.sv:25:5
											VX_elastic_buffer #(
												.DATAW(REQ_DATAW),
												.SIZE(1),
												.OUT_REG(1)
											) req_global_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_valid && is_addr_global),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[282-:4] & ~is_addr_local_mask, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[278], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[277-:120], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[157-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[29-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[13-:12], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[1-:2]}),
												.ready_in(req_global_ready),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].req_valid),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].req_data),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].req_ready)
											);
											// Trace: src/VX_lmem_switch.sv:47:5
											VX_elastic_buffer #(
												.DATAW(REQ_DATAW),
												.SIZE(0),
												.OUT_REG(0)
											) req_local_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_valid && is_addr_local),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[282-:4] & is_addr_local_mask, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[278], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[277-:120], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[157-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[29-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[13-:12], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[1-:2]}),
												.ready_in(req_local_ready),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].req_valid),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].req_data),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].req_ready)
											);
											// Trace: src/VX_lmem_switch.sv:69:5
											VX_stream_arb #(
												.NUM_INPUTS(2),
												.DATAW(RSP_DATAW),
												.ARBITER(ARBITER),
												.OUT_BUF(RSP_OUT_BUF)
											) rsp_arb(
												.clk(clk),
												.reset(reset),
												.valid_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].rsp_valid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].rsp_valid}),
												.ready_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].rsp_ready, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].rsp_ready}),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].rsp_data, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].rsp_data}),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].rsp_data),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].rsp_valid),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].rsp_ready),
												.sel_out()
											);
										end
										assign lmem_switch.clk = clk;
										assign lmem_switch.reset = reset;
									end
									// Trace: src/VX_mem_unit.sv:34:5
									localparam VX_gpu_pkg_LSU_NUM_REQS = 4;
									// expanded interface instance: lmem_bus_if
									localparam _param_4B267_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_4B267_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
									genvar _arr_4B267;
									for (_arr_4B267 = 0; _arr_4B267 <= 3; _arr_4B267 = _arr_4B267 + 1) begin : lmem_bus_if
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_4B267_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_4B267_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_mem_bus_if.sv:7:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_mem_bus_if.sv:9:5
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:21:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire [71:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire [33:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:30:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:31:5
										// Trace: src/VX_mem_bus_if.sv:39:5
									end
									// Trace: src/VX_mem_unit.sv:38:5
									genvar _gv_i_204;
									for (_gv_i_204 = 0; _gv_i_204 < 1; _gv_i_204 = _gv_i_204 + 1) begin : g_lmem_adapters
										localparam i = _gv_i_204;
										// Trace: src/VX_mem_unit.sv:39:9
										// expanded interface instance: lmem_bus_tmp_if
										localparam _param_8C3E5_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
										localparam _param_8C3E5_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
										genvar _arr_8C3E5;
										for (_arr_8C3E5 = 0; _arr_8C3E5 <= 3; _arr_8C3E5 = _arr_8C3E5 + 1) begin : lmem_bus_tmp_if
											// Trace: src/VX_mem_bus_if.sv:2:15
											localparam DATA_SIZE = _param_8C3E5_DATA_SIZE;
											// Trace: src/VX_mem_bus_if.sv:3:15
											localparam FLAGS_WIDTH = 3;
											// Trace: src/VX_mem_bus_if.sv:4:15
											localparam TAG_WIDTH = _param_8C3E5_TAG_WIDTH;
											// Trace: src/VX_mem_bus_if.sv:5:15
											localparam MEM_ADDR_WIDTH = 32;
											// Trace: src/VX_mem_bus_if.sv:6:15
											localparam ADDR_WIDTH = 30;
											// Trace: src/VX_mem_bus_if.sv:7:15
											localparam UUID_WIDTH = 1;
											// Trace: src/VX_mem_bus_if.sv:9:5
											// removed localparam type tag_t
											// Trace: src/VX_mem_bus_if.sv:13:5
											// removed localparam type req_data_t
											// Trace: src/VX_mem_bus_if.sv:21:5
											// removed localparam type rsp_data_t
											// Trace: src/VX_mem_bus_if.sv:25:5
											wire req_valid;
											// Trace: src/VX_mem_bus_if.sv:26:5
											wire [71:0] req_data;
											// Trace: src/VX_mem_bus_if.sv:27:5
											wire req_ready;
											// Trace: src/VX_mem_bus_if.sv:28:5
											wire rsp_valid;
											// Trace: src/VX_mem_bus_if.sv:29:5
											wire [33:0] rsp_data;
											// Trace: src/VX_mem_bus_if.sv:30:5
											wire rsp_ready;
											// Trace: src/VX_mem_bus_if.sv:31:5
											// Trace: src/VX_mem_bus_if.sv:39:5
										end
										// Trace: src/VX_mem_unit.sv:43:9
										// expanded module instance: lmem_adapter
										localparam _bbase_ED918_lsu_mem_if = i;
										localparam _bbase_ED918_mem_bus_if = 0;
										localparam _param_ED918_NUM_LANES = 4;
										localparam _param_ED918_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
										localparam _param_ED918_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
										localparam _param_ED918_TAG_SEL_BITS = 1;
										localparam _param_ED918_ARBITER = "P";
										localparam _param_ED918_REQ_OUT_BUF = 3;
										localparam _param_ED918_RSP_OUT_BUF = 2;
										if (1) begin : lmem_adapter
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_lsu_adapter.sv:2:15
											localparam NUM_LANES = _param_ED918_NUM_LANES;
											// Trace: src/VX_lsu_adapter.sv:3:15
											localparam DATA_SIZE = _param_ED918_DATA_SIZE;
											// Trace: src/VX_lsu_adapter.sv:4:15
											localparam TAG_WIDTH = _param_ED918_TAG_WIDTH;
											// Trace: src/VX_lsu_adapter.sv:5:15
											localparam TAG_SEL_BITS = _param_ED918_TAG_SEL_BITS;
											// Trace: src/VX_lsu_adapter.sv:6:16
											localparam ARBITER = _param_ED918_ARBITER;
											// Trace: src/VX_lsu_adapter.sv:7:15
											localparam REQ_OUT_BUF = _param_ED918_REQ_OUT_BUF;
											// Trace: src/VX_lsu_adapter.sv:8:15
											localparam RSP_OUT_BUF = _param_ED918_RSP_OUT_BUF;
											// Trace: src/VX_lsu_adapter.sv:10:5
											wire clk;
											// Trace: src/VX_lsu_adapter.sv:11:5
											wire reset;
											// Trace: src/VX_lsu_adapter.sv:12:5
											localparam _mbase_lsu_mem_if = _bbase_ED918_lsu_mem_if;
											// Trace: src/VX_lsu_adapter.sv:13:5
											localparam _mbase_mem_bus_if = 0;
											// Trace: src/VX_lsu_adapter.sv:15:5
											localparam REQ_ADDR_WIDTH = 30;
											// Trace: src/VX_lsu_adapter.sv:16:5
											localparam REQ_DATA_WIDTH = 70;
											// Trace: src/VX_lsu_adapter.sv:17:5
											localparam RSP_DATA_WIDTH = 32;
											// Trace: src/VX_lsu_adapter.sv:18:5
											wire [279:0] req_data_in;
											// Trace: src/VX_lsu_adapter.sv:19:5
											wire [3:0] req_valid_out;
											// Trace: src/VX_lsu_adapter.sv:20:5
											wire [279:0] req_data_out;
											// Trace: src/VX_lsu_adapter.sv:21:5
											wire [7:0] req_tag_out;
											// Trace: src/VX_lsu_adapter.sv:22:5
											wire [3:0] req_ready_out;
											// Trace: src/VX_lsu_adapter.sv:23:5
											genvar _gv_i_148;
											for (_gv_i_148 = 0; _gv_i_148 < NUM_LANES; _gv_i_148 = _gv_i_148 + 1) begin : g_req_data_in
												localparam i = _gv_i_148;
												// Trace: src/VX_lsu_adapter.sv:24:9
												assign req_data_in[i * 70+:70] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].req_data[278], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].req_data[158 + (i * 30)+:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].req_data[30 + (i * 32)+:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].req_data[14 + (i * 4)+:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].req_data[2 + (i * 3)+:3]};
											end
											// Trace: src/VX_lsu_adapter.sv:32:5
											VX_stream_unpack #(
												.NUM_REQS(NUM_LANES),
												.DATA_WIDTH(REQ_DATA_WIDTH),
												.TAG_WIDTH(TAG_WIDTH),
												.OUT_BUF(REQ_OUT_BUF)
											) stream_unpack(
												.clk(clk),
												.reset(reset),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].req_valid),
												.mask_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].req_data[282-:4]),
												.data_in(req_data_in),
												.tag_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].req_data[1-:2]),
												.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].req_ready),
												.valid_out(req_valid_out),
												.data_out(req_data_out),
												.tag_out(req_tag_out),
												.ready_out(req_ready_out)
											);
											// Trace: src/VX_lsu_adapter.sv:50:5
											genvar _gv_i_149;
											for (_gv_i_149 = 0; _gv_i_149 < NUM_LANES; _gv_i_149 = _gv_i_149 + 1) begin : g_mem_bus_req
												localparam i = _gv_i_149;
												// Trace: src/VX_lsu_adapter.sv:51:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].req_valid = req_valid_out[i];
												// Trace: src/VX_lsu_adapter.sv:52:9
												assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].req_data[71], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].req_data[70-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].req_data[40-:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].req_data[8-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].req_data[4-:3]} = req_data_out[i * 70+:70];
												// Trace: src/VX_lsu_adapter.sv:59:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].req_data[1-:2] = req_tag_out[i * 2+:2];
												// Trace: src/VX_lsu_adapter.sv:60:9
												assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].req_ready;
											end
											// Trace: src/VX_lsu_adapter.sv:62:5
											wire [3:0] rsp_valid_out;
											// Trace: src/VX_lsu_adapter.sv:63:5
											wire [127:0] rsp_data_out;
											// Trace: src/VX_lsu_adapter.sv:64:5
											wire [7:0] rsp_tag_out;
											// Trace: src/VX_lsu_adapter.sv:65:5
											wire [3:0] rsp_ready_out;
											// Trace: src/VX_lsu_adapter.sv:66:5
											genvar _gv_i_150;
											for (_gv_i_150 = 0; _gv_i_150 < NUM_LANES; _gv_i_150 = _gv_i_150 + 1) begin : g_mem_bus_rsp
												localparam i = _gv_i_150;
												// Trace: src/VX_lsu_adapter.sv:67:9
												assign rsp_valid_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].rsp_valid;
												// Trace: src/VX_lsu_adapter.sv:68:9
												assign rsp_data_out[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].rsp_data[33-:32];
												// Trace: src/VX_lsu_adapter.sv:69:9
												assign rsp_tag_out[i * 2+:2] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].rsp_data[1-:2];
												// Trace: src/VX_lsu_adapter.sv:70:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_lmem_adapters[_gv_i_204].lmem_bus_tmp_if[i + _mbase_mem_bus_if].rsp_ready = rsp_ready_out[i];
											end
											// Trace: src/VX_lsu_adapter.sv:72:5
											VX_stream_pack #(
												.NUM_REQS(NUM_LANES),
												.DATA_WIDTH(RSP_DATA_WIDTH),
												.TAG_WIDTH(TAG_WIDTH),
												.TAG_SEL_BITS(TAG_SEL_BITS),
												.ARBITER(ARBITER),
												.OUT_BUF(RSP_OUT_BUF)
											) stream_pack(
												.clk(clk),
												.reset(reset),
												.valid_in(rsp_valid_out),
												.data_in(rsp_data_out),
												.tag_in(rsp_tag_out),
												.ready_in(rsp_ready_out),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].rsp_valid),
												.mask_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].rsp_data[133-:4]),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].rsp_data[129-:128]),
												.tag_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].rsp_data[1-:2]),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_lsu_mem_if].rsp_ready)
											);
										end
										assign lmem_adapter.clk = clk;
										assign lmem_adapter.reset = reset;
										genvar _gv_j_20;
										for (_gv_j_20 = 0; _gv_j_20 < 4; _gv_j_20 = _gv_j_20 + 1) begin : g_lmem_bus_if
											localparam j = _gv_j_20;
											// Trace: src/VX_mem_unit.sv:58:5
											assign lmem_bus_if[(i * 4) + j].req_valid = lmem_bus_tmp_if[j].req_valid;
											// Trace: src/VX_mem_unit.sv:59:5
											assign lmem_bus_if[(i * 4) + j].req_data = lmem_bus_tmp_if[j].req_data;
											// Trace: src/VX_mem_unit.sv:60:5
											assign lmem_bus_tmp_if[j].req_ready = lmem_bus_if[(i * 4) + j].req_ready;
											// Trace: src/VX_mem_unit.sv:61:5
											assign lmem_bus_tmp_if[j].rsp_valid = lmem_bus_if[(i * 4) + j].rsp_valid;
											// Trace: src/VX_mem_unit.sv:62:5
											assign lmem_bus_tmp_if[j].rsp_data = lmem_bus_if[(i * 4) + j].rsp_data;
											// Trace: src/VX_mem_unit.sv:63:5
											assign lmem_bus_if[(i * 4) + j].rsp_ready = lmem_bus_tmp_if[j].rsp_ready;
										end
									end
									// Trace: src/VX_mem_unit.sv:66:5
									// expanded module instance: local_mem
									localparam _bbase_9EDEE_mem_bus_if = 0;
									localparam _param_9EDEE_INSTANCE_ID = "";
									localparam _param_9EDEE_SIZE = 16384;
									localparam _param_9EDEE_NUM_REQS = VX_gpu_pkg_LSU_NUM_REQS;
									localparam _param_9EDEE_NUM_BANKS = 4;
									localparam _param_9EDEE_WORD_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_9EDEE_ADDR_WIDTH = LMEM_ADDR_WIDTH;
									localparam _param_9EDEE_UUID_WIDTH = 1;
									localparam _param_9EDEE_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
									localparam _param_9EDEE_OUT_BUF = 3;
									if (1) begin : local_mem
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_local_mem.sv:2:17
										localparam INSTANCE_ID = _param_9EDEE_INSTANCE_ID;
										// Trace: src/VX_local_mem.sv:3:15
										localparam SIZE = _param_9EDEE_SIZE;
										// Trace: src/VX_local_mem.sv:4:15
										localparam NUM_REQS = _param_9EDEE_NUM_REQS;
										// Trace: src/VX_local_mem.sv:5:15
										localparam NUM_BANKS = _param_9EDEE_NUM_BANKS;
										// Trace: src/VX_local_mem.sv:6:15
										localparam ADDR_WIDTH = _param_9EDEE_ADDR_WIDTH;
										// Trace: src/VX_local_mem.sv:7:15
										localparam WORD_SIZE = _param_9EDEE_WORD_SIZE;
										// Trace: src/VX_local_mem.sv:8:15
										localparam UUID_WIDTH = _param_9EDEE_UUID_WIDTH;
										// Trace: src/VX_local_mem.sv:9:15
										localparam TAG_WIDTH = _param_9EDEE_TAG_WIDTH;
										// Trace: src/VX_local_mem.sv:10:15
										localparam OUT_BUF = _param_9EDEE_OUT_BUF;
										// Trace: src/VX_local_mem.sv:12:5
										wire clk;
										// Trace: src/VX_local_mem.sv:13:5
										wire reset;
										// Trace: src/VX_local_mem.sv:14:5
										localparam _mbase_mem_bus_if = 0;
										// Trace: src/VX_local_mem.sv:16:5
										localparam REQ_SEL_BITS = 2;
										// Trace: src/VX_local_mem.sv:17:5
										localparam REQ_SEL_WIDTH = REQ_SEL_BITS;
										// Trace: src/VX_local_mem.sv:18:5
										localparam WORD_WIDTH = 32;
										// Trace: src/VX_local_mem.sv:19:5
										localparam NUM_WORDS = 4096;
										// Trace: src/VX_local_mem.sv:20:5
										localparam WORDS_PER_BANK = 1024;
										// Trace: src/VX_local_mem.sv:21:5
										localparam BANK_ADDR_WIDTH = 10;
										// Trace: src/VX_local_mem.sv:22:5
										localparam BANK_SEL_BITS = 2;
										// Trace: src/VX_local_mem.sv:23:5
										localparam BANK_SEL_WIDTH = BANK_SEL_BITS;
										// Trace: src/VX_local_mem.sv:24:5
										localparam REQ_DATAW = 49;
										// Trace: src/VX_local_mem.sv:25:5
										localparam RSP_DATAW = 34;
										// Trace: src/VX_local_mem.sv:26:5
										wire [7:0] req_bank_idx;
										// Trace: src/VX_local_mem.sv:27:5
										if (1) begin : g_req_bank_idx
											genvar _gv_i_72;
											for (_gv_i_72 = 0; _gv_i_72 < NUM_REQS; _gv_i_72 = _gv_i_72 + 1) begin : g_req_bank_idxs
												localparam i = _gv_i_72;
												// Trace: src/VX_local_mem.sv:29:13
												assign req_bank_idx[i * 2+:2] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].req_data[41+:BANK_SEL_BITS];
											end
										end
										// Trace: src/VX_local_mem.sv:34:5
										wire [39:0] req_bank_addr;
										// Trace: src/VX_local_mem.sv:35:5
										genvar _gv_i_73;
										for (_gv_i_73 = 0; _gv_i_73 < NUM_REQS; _gv_i_73 = _gv_i_73 + 1) begin : g_req_bank_addr
											localparam i = _gv_i_73;
											// Trace: src/VX_local_mem.sv:36:9
											assign req_bank_addr[i * 10+:10] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].req_data[43+:BANK_ADDR_WIDTH];
										end
										// Trace: src/VX_local_mem.sv:38:5
										wire [3:0] per_bank_req_valid;
										// Trace: src/VX_local_mem.sv:39:5
										wire [3:0] per_bank_req_rw;
										// Trace: src/VX_local_mem.sv:40:5
										wire [39:0] per_bank_req_addr;
										// Trace: src/VX_local_mem.sv:41:5
										wire [15:0] per_bank_req_byteen;
										// Trace: src/VX_local_mem.sv:42:5
										wire [127:0] per_bank_req_data;
										// Trace: src/VX_local_mem.sv:43:5
										wire [7:0] per_bank_req_tag;
										// Trace: src/VX_local_mem.sv:44:5
										wire [7:0] per_bank_req_idx;
										// Trace: src/VX_local_mem.sv:45:5
										wire [3:0] per_bank_req_ready;
										// Trace: src/VX_local_mem.sv:46:5
										wire [195:0] per_bank_req_data_aos;
										// Trace: src/VX_local_mem.sv:47:5
										wire [3:0] req_valid_in;
										// Trace: src/VX_local_mem.sv:48:5
										wire [195:0] req_data_in;
										// Trace: src/VX_local_mem.sv:49:5
										wire [3:0] req_ready_in;
										// Trace: src/VX_local_mem.sv:50:5
										genvar _gv_i_74;
										for (_gv_i_74 = 0; _gv_i_74 < NUM_REQS; _gv_i_74 = _gv_i_74 + 1) begin : g_req_data_in
											localparam i = _gv_i_74;
											// Trace: src/VX_local_mem.sv:51:9
											assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].req_valid;
											// Trace: src/VX_local_mem.sv:52:9
											assign req_data_in[i * 49+:49] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].req_data[71], req_bank_addr[i * 10+:10], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].req_data[40-:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].req_data[8-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].req_data[1-:2]};
											// Trace: src/VX_local_mem.sv:59:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].req_ready = req_ready_in[i];
										end
										// Trace: src/VX_local_mem.sv:61:5
										VX_stream_xbar #(
											.NUM_INPUTS(NUM_REQS),
											.NUM_OUTPUTS(NUM_BANKS),
											.DATAW(REQ_DATAW),
											.PERF_CTR_BITS(44),
											.ARBITER("P"),
											.OUT_BUF(3)
										) req_xbar(
											.clk(clk),
											.reset(reset),
											.collisions(),
											.valid_in(req_valid_in),
											.data_in(req_data_in),
											.sel_in(req_bank_idx),
											.ready_in(req_ready_in),
											.valid_out(per_bank_req_valid),
											.data_out(per_bank_req_data_aos),
											.sel_out(per_bank_req_idx),
											.ready_out(per_bank_req_ready)
										);
										// Trace: src/VX_local_mem.sv:81:5
										genvar _gv_i_75;
										for (_gv_i_75 = 0; _gv_i_75 < NUM_BANKS; _gv_i_75 = _gv_i_75 + 1) begin : g_per_bank_req_data_soa
											localparam i = _gv_i_75;
											// Trace: src/VX_local_mem.sv:82:9
											assign {per_bank_req_rw[i], per_bank_req_addr[i * 10+:10], per_bank_req_data[i * 32+:32], per_bank_req_byteen[i * 4+:4], per_bank_req_tag[i * 2+:2]} = per_bank_req_data_aos[i * 49+:49];
										end
										// Trace: src/VX_local_mem.sv:90:5
										wire [3:0] per_bank_rsp_valid;
										// Trace: src/VX_local_mem.sv:91:5
										wire [127:0] per_bank_rsp_data;
										// Trace: src/VX_local_mem.sv:92:5
										wire [7:0] per_bank_rsp_idx;
										// Trace: src/VX_local_mem.sv:93:5
										wire [7:0] per_bank_rsp_tag;
										// Trace: src/VX_local_mem.sv:94:5
										wire [3:0] per_bank_rsp_ready;
										// Trace: src/VX_local_mem.sv:95:5
										genvar _gv_i_76;
										for (_gv_i_76 = 0; _gv_i_76 < NUM_BANKS; _gv_i_76 = _gv_i_76 + 1) begin : g_data_store
											localparam i = _gv_i_76;
											// Trace: src/VX_local_mem.sv:96:9
											wire bank_rsp_valid;
											wire bank_rsp_ready;
											// Trace: src/VX_local_mem.sv:97:9
											VX_sp_ram #(
												.DATAW(WORD_WIDTH),
												.SIZE(WORDS_PER_BANK),
												.WRENW(WORD_SIZE),
												.OUT_REG(1),
												.RDW_MODE("R")
											) lmem_store(
												.clk(clk),
												.reset(reset),
												.read((per_bank_req_valid[i] && per_bank_req_ready[i]) && ~per_bank_req_rw[i]),
												.write((per_bank_req_valid[i] && per_bank_req_ready[i]) && per_bank_req_rw[i]),
												.wren(per_bank_req_byteen[i * 4+:4]),
												.addr(per_bank_req_addr[i * 10+:10]),
												.wdata(per_bank_req_data[i * 32+:32]),
												.rdata(per_bank_rsp_data[i * 32+:32])
											);
											// Trace: src/VX_local_mem.sv:113:9
											reg [9:0] last_wr_addr;
											// Trace: src/VX_local_mem.sv:114:9
											reg last_wr_valid;
											// Trace: src/VX_local_mem.sv:115:9
											always @(posedge clk) begin
												// Trace: src/VX_local_mem.sv:116:13
												if (reset)
													// Trace: src/VX_local_mem.sv:117:17
													last_wr_valid <= 0;
												else
													// Trace: src/VX_local_mem.sv:119:17
													last_wr_valid <= (per_bank_req_valid[i] && per_bank_req_ready[i]) && per_bank_req_rw[i];
												// Trace: src/VX_local_mem.sv:121:13
												last_wr_addr <= per_bank_req_addr[i * 10+:10];
											end
											// Trace: src/VX_local_mem.sv:123:9
											wire is_rdw_hazard = (last_wr_valid && ~per_bank_req_rw[i]) && (per_bank_req_addr[i * 10+:10] == last_wr_addr);
											// Trace: src/VX_local_mem.sv:124:9
											assign bank_rsp_valid = (per_bank_req_valid[i] && ~per_bank_req_rw[i]) && ~is_rdw_hazard;
											// Trace: src/VX_local_mem.sv:125:9
											assign per_bank_req_ready[i] = (bank_rsp_ready || per_bank_req_rw[i]) && ~is_rdw_hazard;
											// Trace: src/VX_local_mem.sv:126:9
											VX_pipe_buffer #(.DATAW(4)) bram_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(bank_rsp_valid),
												.ready_in(bank_rsp_ready),
												.data_in({per_bank_req_idx[i * 2+:2], per_bank_req_tag[i * 2+:2]}),
												.data_out({per_bank_rsp_idx[i * 2+:2], per_bank_rsp_tag[i * 2+:2]}),
												.valid_out(per_bank_rsp_valid[i]),
												.ready_out(per_bank_rsp_ready[i])
											);
										end
										// Trace: src/VX_local_mem.sv:139:5
										wire [135:0] per_bank_rsp_data_aos;
										// Trace: src/VX_local_mem.sv:140:5
										genvar _gv_i_77;
										for (_gv_i_77 = 0; _gv_i_77 < NUM_BANKS; _gv_i_77 = _gv_i_77 + 1) begin : g_per_bank_rsp_data_aos
											localparam i = _gv_i_77;
											// Trace: src/VX_local_mem.sv:141:9
											assign per_bank_rsp_data_aos[i * 34+:34] = {per_bank_rsp_data[i * 32+:32], per_bank_rsp_tag[i * 2+:2]};
										end
										// Trace: src/VX_local_mem.sv:143:5
										wire [3:0] rsp_valid_out;
										// Trace: src/VX_local_mem.sv:144:5
										wire [135:0] rsp_data_out;
										// Trace: src/VX_local_mem.sv:145:5
										wire [3:0] rsp_ready_out;
										// Trace: src/VX_local_mem.sv:146:5
										VX_stream_xbar #(
											.NUM_INPUTS(NUM_BANKS),
											.NUM_OUTPUTS(NUM_REQS),
											.DATAW(RSP_DATAW),
											.ARBITER("P"),
											.OUT_BUF(OUT_BUF)
										) rsp_xbar(
											.clk(clk),
											.reset(reset),
											.collisions(),
											.sel_in(per_bank_rsp_idx),
											.valid_in(per_bank_rsp_valid),
											.data_in(per_bank_rsp_data_aos),
											.ready_in(per_bank_rsp_ready),
											.valid_out(rsp_valid_out),
											.data_out(rsp_data_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
										// Trace: src/VX_local_mem.sv:165:5
										genvar _gv_i_78;
										for (_gv_i_78 = 0; _gv_i_78 < NUM_REQS; _gv_i_78 = _gv_i_78 + 1) begin : g_mem_bus_if
											localparam i = _gv_i_78;
											// Trace: src/VX_local_mem.sv:166:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].rsp_valid = rsp_valid_out[i];
											// Trace: src/VX_local_mem.sv:167:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].rsp_data = rsp_data_out[i * 34+:34];
											// Trace: src/VX_local_mem.sv:168:9
											assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_bus_if[i + _mbase_mem_bus_if].rsp_ready;
										end
									end
									assign local_mem.clk = clk;
									assign local_mem.reset = reset;
									// Trace: src/VX_mem_unit.sv:81:5
									localparam VX_gpu_pkg_DCACHE_MERGED_REQS = 1;
									localparam VX_gpu_pkg_DCACHE_MEM_BATCHES = 1;
									localparam VX_gpu_pkg_DCACHE_TAG_ID_BITS = 2;
									localparam VX_gpu_pkg_DCACHE_TAG_WIDTH = 3;
									// expanded interface instance: dcache_coalesced_if
									localparam _param_419A9_NUM_LANES = VX_gpu_pkg_DCACHE_CHANNELS;
									localparam _param_419A9_DATA_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
									localparam _param_419A9_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
									genvar _arr_419A9;
									for (_arr_419A9 = 0; _arr_419A9 <= 0; _arr_419A9 = _arr_419A9 + 1) begin : dcache_coalesced_if
										// Trace: src/VX_lsu_mem_if.sv:2:15
										localparam NUM_LANES = _param_419A9_NUM_LANES;
										// Trace: src/VX_lsu_mem_if.sv:3:15
										localparam DATA_SIZE = _param_419A9_DATA_SIZE;
										// Trace: src/VX_lsu_mem_if.sv:4:15
										localparam TAG_WIDTH = _param_419A9_TAG_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:5:15
										localparam FLAGS_WIDTH = 3;
										// Trace: src/VX_lsu_mem_if.sv:6:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_lsu_mem_if.sv:7:15
										localparam ADDR_WIDTH = 28;
										// Trace: src/VX_lsu_mem_if.sv:8:15
										localparam UUID_WIDTH = 1;
										// Trace: src/VX_lsu_mem_if.sv:10:5
										// removed localparam type tag_t
										// Trace: src/VX_lsu_mem_if.sv:14:5
										// removed localparam type req_data_t
										// Trace: src/VX_lsu_mem_if.sv:23:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_lsu_mem_if.sv:28:5
										wire req_valid;
										// Trace: src/VX_lsu_mem_if.sv:29:5
										wire [179:0] req_data;
										// Trace: src/VX_lsu_mem_if.sv:30:5
										wire req_ready;
										// Trace: src/VX_lsu_mem_if.sv:31:5
										wire rsp_valid;
										// Trace: src/VX_lsu_mem_if.sv:32:5
										wire [131:0] rsp_data;
										// Trace: src/VX_lsu_mem_if.sv:33:5
										wire rsp_ready;
										// Trace: src/VX_lsu_mem_if.sv:34:5
										// Trace: src/VX_lsu_mem_if.sv:42:5
									end
									// Trace: src/VX_mem_unit.sv:86:5
									localparam VX_gpu_pkg_LSU_ADDR_WIDTH = 30;
									if (1) begin : g_enabled
										genvar _gv_i_205;
										for (_gv_i_205 = 0; _gv_i_205 < 1; _gv_i_205 = _gv_i_205 + 1) begin : g_coalescers
											localparam i = _gv_i_205;
											// Trace: src/VX_mem_unit.sv:88:13
											VX_mem_coalescer #(
												.INSTANCE_ID(""),
												.NUM_REQS(4),
												.DATA_IN_SIZE(VX_gpu_pkg_LSU_WORD_SIZE),
												.DATA_OUT_SIZE(VX_gpu_pkg_DCACHE_WORD_SIZE),
												.ADDR_WIDTH(VX_gpu_pkg_LSU_ADDR_WIDTH),
												.FLAGS_WIDTH(3),
												.TAG_WIDTH(VX_gpu_pkg_LSU_TAG_WIDTH),
												.UUID_WIDTH(1),
												.QUEUE_SIZE(4)
											) mem_coalescer(
												.clk(clk),
												.reset(reset),
												.in_req_valid(lsu_dcache_if[i].req_valid),
												.in_req_mask(lsu_dcache_if[i].req_data[282-:4]),
												.in_req_rw(lsu_dcache_if[i].req_data[278]),
												.in_req_byteen(lsu_dcache_if[i].req_data[29-:16]),
												.in_req_addr(lsu_dcache_if[i].req_data[277-:120]),
												.in_req_flags(lsu_dcache_if[i].req_data[13-:12]),
												.in_req_data(lsu_dcache_if[i].req_data[157-:128]),
												.in_req_tag(lsu_dcache_if[i].req_data[1-:2]),
												.in_req_ready(lsu_dcache_if[i].req_ready),
												.in_rsp_valid(lsu_dcache_if[i].rsp_valid),
												.in_rsp_mask(lsu_dcache_if[i].rsp_data[133-:4]),
												.in_rsp_data(lsu_dcache_if[i].rsp_data[129-:128]),
												.in_rsp_tag(lsu_dcache_if[i].rsp_data[1-:2]),
												.in_rsp_ready(lsu_dcache_if[i].rsp_ready),
												.out_req_valid(dcache_coalesced_if[i].req_valid),
												.out_req_mask(dcache_coalesced_if[i].req_data[179-:1]),
												.out_req_rw(dcache_coalesced_if[i].req_data[178]),
												.out_req_byteen(dcache_coalesced_if[i].req_data[21-:16]),
												.out_req_addr(dcache_coalesced_if[i].req_data[177-:28]),
												.out_req_flags(dcache_coalesced_if[i].req_data[5-:3]),
												.out_req_data(dcache_coalesced_if[i].req_data[149-:128]),
												.out_req_tag(dcache_coalesced_if[i].req_data[2-:3]),
												.out_req_ready(dcache_coalesced_if[i].req_ready),
												.out_rsp_valid(dcache_coalesced_if[i].rsp_valid),
												.out_rsp_mask(dcache_coalesced_if[i].rsp_data[131-:1]),
												.out_rsp_data(dcache_coalesced_if[i].rsp_data[130-:128]),
												.out_rsp_tag(dcache_coalesced_if[i].rsp_data[2-:3]),
												.out_rsp_ready(dcache_coalesced_if[i].rsp_ready)
											);
										end
									end
									// Trace: src/VX_mem_unit.sv:141:5
									genvar _gv_i_207;
									for (_gv_i_207 = 0; _gv_i_207 < 1; _gv_i_207 = _gv_i_207 + 1) begin : g_dcache_adapters
										localparam i = _gv_i_207;
										// Trace: src/VX_mem_unit.sv:142:9
										// expanded interface instance: dcache_bus_tmp_if
										localparam _param_CE5A6_DATA_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
										localparam _param_CE5A6_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
										genvar _arr_CE5A6;
										for (_arr_CE5A6 = 0; _arr_CE5A6 <= 0; _arr_CE5A6 = _arr_CE5A6 + 1) begin : dcache_bus_tmp_if
											// Trace: src/VX_mem_bus_if.sv:2:15
											localparam DATA_SIZE = _param_CE5A6_DATA_SIZE;
											// Trace: src/VX_mem_bus_if.sv:3:15
											localparam FLAGS_WIDTH = 3;
											// Trace: src/VX_mem_bus_if.sv:4:15
											localparam TAG_WIDTH = _param_CE5A6_TAG_WIDTH;
											// Trace: src/VX_mem_bus_if.sv:5:15
											localparam MEM_ADDR_WIDTH = 32;
											// Trace: src/VX_mem_bus_if.sv:6:15
											localparam ADDR_WIDTH = 28;
											// Trace: src/VX_mem_bus_if.sv:7:15
											localparam UUID_WIDTH = 1;
											// Trace: src/VX_mem_bus_if.sv:9:5
											// removed localparam type tag_t
											// Trace: src/VX_mem_bus_if.sv:13:5
											// removed localparam type req_data_t
											// Trace: src/VX_mem_bus_if.sv:21:5
											// removed localparam type rsp_data_t
											// Trace: src/VX_mem_bus_if.sv:25:5
											wire req_valid;
											// Trace: src/VX_mem_bus_if.sv:26:5
											wire [178:0] req_data;
											// Trace: src/VX_mem_bus_if.sv:27:5
											wire req_ready;
											// Trace: src/VX_mem_bus_if.sv:28:5
											wire rsp_valid;
											// Trace: src/VX_mem_bus_if.sv:29:5
											wire [130:0] rsp_data;
											// Trace: src/VX_mem_bus_if.sv:30:5
											wire rsp_ready;
											// Trace: src/VX_mem_bus_if.sv:31:5
											// Trace: src/VX_mem_bus_if.sv:39:5
										end
										// Trace: src/VX_mem_unit.sv:146:9
										// expanded module instance: dcache_adapter
										localparam _bbase_6EE01_lsu_mem_if = i;
										localparam _bbase_6EE01_mem_bus_if = 0;
										localparam _param_6EE01_NUM_LANES = VX_gpu_pkg_DCACHE_CHANNELS;
										localparam _param_6EE01_DATA_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
										localparam _param_6EE01_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
										localparam _param_6EE01_TAG_SEL_BITS = 2;
										localparam _param_6EE01_ARBITER = "P";
										localparam _param_6EE01_REQ_OUT_BUF = 0;
										localparam _param_6EE01_RSP_OUT_BUF = 0;
										if (1) begin : dcache_adapter
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_lsu_adapter.sv:2:15
											localparam NUM_LANES = _param_6EE01_NUM_LANES;
											// Trace: src/VX_lsu_adapter.sv:3:15
											localparam DATA_SIZE = _param_6EE01_DATA_SIZE;
											// Trace: src/VX_lsu_adapter.sv:4:15
											localparam TAG_WIDTH = _param_6EE01_TAG_WIDTH;
											// Trace: src/VX_lsu_adapter.sv:5:15
											localparam TAG_SEL_BITS = _param_6EE01_TAG_SEL_BITS;
											// Trace: src/VX_lsu_adapter.sv:6:16
											localparam ARBITER = _param_6EE01_ARBITER;
											// Trace: src/VX_lsu_adapter.sv:7:15
											localparam REQ_OUT_BUF = _param_6EE01_REQ_OUT_BUF;
											// Trace: src/VX_lsu_adapter.sv:8:15
											localparam RSP_OUT_BUF = _param_6EE01_RSP_OUT_BUF;
											// Trace: src/VX_lsu_adapter.sv:10:5
											wire clk;
											// Trace: src/VX_lsu_adapter.sv:11:5
											wire reset;
											// Trace: src/VX_lsu_adapter.sv:12:5
											localparam _mbase_lsu_mem_if = _bbase_6EE01_lsu_mem_if;
											// Trace: src/VX_lsu_adapter.sv:13:5
											localparam _mbase_mem_bus_if = 0;
											// Trace: src/VX_lsu_adapter.sv:15:5
											localparam REQ_ADDR_WIDTH = 28;
											// Trace: src/VX_lsu_adapter.sv:16:5
											localparam REQ_DATA_WIDTH = 176;
											// Trace: src/VX_lsu_adapter.sv:17:5
											localparam RSP_DATA_WIDTH = 128;
											// Trace: src/VX_lsu_adapter.sv:18:5
											wire [175:0] req_data_in;
											// Trace: src/VX_lsu_adapter.sv:19:5
											wire [0:0] req_valid_out;
											// Trace: src/VX_lsu_adapter.sv:20:5
											wire [175:0] req_data_out;
											// Trace: src/VX_lsu_adapter.sv:21:5
											wire [2:0] req_tag_out;
											// Trace: src/VX_lsu_adapter.sv:22:5
											wire [0:0] req_ready_out;
											// Trace: src/VX_lsu_adapter.sv:23:5
											genvar _gv_i_148;
											for (_gv_i_148 = 0; _gv_i_148 < NUM_LANES; _gv_i_148 = _gv_i_148 + 1) begin : g_req_data_in
												localparam i = _gv_i_148;
												// Trace: src/VX_lsu_adapter.sv:24:9
												assign req_data_in[i * 176+:176] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[178], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[150 + (i * 28)+:28], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[22 + (i * 128)+:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[6 + (i * 16)+:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[3 + (i * 3)+:3]};
											end
											// Trace: src/VX_lsu_adapter.sv:32:5
											VX_stream_unpack #(
												.NUM_REQS(NUM_LANES),
												.DATA_WIDTH(REQ_DATA_WIDTH),
												.TAG_WIDTH(TAG_WIDTH),
												.OUT_BUF(REQ_OUT_BUF)
											) stream_unpack(
												.clk(clk),
												.reset(reset),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_valid),
												.mask_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[179-:1]),
												.data_in(req_data_in),
												.tag_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[2-:3]),
												.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_ready),
												.valid_out(req_valid_out),
												.data_out(req_data_out),
												.tag_out(req_tag_out),
												.ready_out(req_ready_out)
											);
											// Trace: src/VX_lsu_adapter.sv:50:5
											genvar _gv_i_149;
											for (_gv_i_149 = 0; _gv_i_149 < NUM_LANES; _gv_i_149 = _gv_i_149 + 1) begin : g_mem_bus_req
												localparam i = _gv_i_149;
												// Trace: src/VX_lsu_adapter.sv:51:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_valid = req_valid_out[i];
												// Trace: src/VX_lsu_adapter.sv:52:9
												assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[178], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[177-:28], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[149-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[21-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[5-:3]} = req_data_out[i * 176+:176];
												// Trace: src/VX_lsu_adapter.sv:59:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[2-:3] = req_tag_out[i * 3+:3];
												// Trace: src/VX_lsu_adapter.sv:60:9
												assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_ready;
											end
											// Trace: src/VX_lsu_adapter.sv:62:5
											wire [0:0] rsp_valid_out;
											// Trace: src/VX_lsu_adapter.sv:63:5
											wire [127:0] rsp_data_out;
											// Trace: src/VX_lsu_adapter.sv:64:5
											wire [2:0] rsp_tag_out;
											// Trace: src/VX_lsu_adapter.sv:65:5
											wire [0:0] rsp_ready_out;
											// Trace: src/VX_lsu_adapter.sv:66:5
											genvar _gv_i_150;
											for (_gv_i_150 = 0; _gv_i_150 < NUM_LANES; _gv_i_150 = _gv_i_150 + 1) begin : g_mem_bus_rsp
												localparam i = _gv_i_150;
												// Trace: src/VX_lsu_adapter.sv:67:9
												assign rsp_valid_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].rsp_valid;
												// Trace: src/VX_lsu_adapter.sv:68:9
												assign rsp_data_out[i * 128+:128] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].rsp_data[130-:128];
												// Trace: src/VX_lsu_adapter.sv:69:9
												assign rsp_tag_out[i * 3+:3] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].rsp_data[2-:3];
												// Trace: src/VX_lsu_adapter.sv:70:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_207].dcache_bus_tmp_if[i + _mbase_mem_bus_if].rsp_ready = rsp_ready_out[i];
											end
											// Trace: src/VX_lsu_adapter.sv:72:5
											VX_stream_pack #(
												.NUM_REQS(NUM_LANES),
												.DATA_WIDTH(RSP_DATA_WIDTH),
												.TAG_WIDTH(TAG_WIDTH),
												.TAG_SEL_BITS(TAG_SEL_BITS),
												.ARBITER(ARBITER),
												.OUT_BUF(RSP_OUT_BUF)
											) stream_pack(
												.clk(clk),
												.reset(reset),
												.valid_in(rsp_valid_out),
												.data_in(rsp_data_out),
												.tag_in(rsp_tag_out),
												.ready_in(rsp_ready_out),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_valid),
												.mask_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_data[131-:1]),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_data[130-:128]),
												.tag_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_data[2-:3]),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_ready)
											);
										end
										assign dcache_adapter.clk = clk;
										assign dcache_adapter.reset = reset;
										genvar _gv_j_21;
										for (_gv_j_21 = 0; _gv_j_21 < VX_gpu_pkg_DCACHE_CHANNELS; _gv_j_21 = _gv_j_21 + 1) begin : g_dcache_bus_if
											localparam j = _gv_j_21;
											// Trace: src/VX_mem_unit.sv:161:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].req_valid = dcache_bus_tmp_if[j].req_valid;
											// Trace: src/VX_mem_unit.sv:162:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].req_data = dcache_bus_tmp_if[j].req_data;
											// Trace: src/VX_mem_unit.sv:163:5
											assign dcache_bus_tmp_if[j].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].req_ready;
											// Trace: src/VX_mem_unit.sv:164:5
											assign dcache_bus_tmp_if[j].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].rsp_valid;
											// Trace: src/VX_mem_unit.sv:165:5
											assign dcache_bus_tmp_if[j].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].rsp_data;
											// Trace: src/VX_mem_unit.sv:166:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].rsp_ready = dcache_bus_tmp_if[j].rsp_ready;
										end
									end
								end
								assign mem_unit.clk = clk;
								assign mem_unit.reset = reset;
							end
							assign core.clk = clk;
							assign core.reset = core_reset;
							assign per_core_busy[core_id] = core.busy;
						end
						// Trace: src/VX_socket.sv:325:5
						VX_pipe_register #(
							.DATAW(1),
							.RESETW(1),
							.DEPTH(1'd0)
						) __busy__(
							.clk(clk),
							.reset(reset),
							.enable(1'b1),
							.data_in(|per_core_busy),
							.data_out(busy)
						);
					end
					assign socket.clk = clk;
					assign socket.reset = socket_reset;
					assign per_socket_busy[socket_id] = socket.busy;
				end
				// Trace: src/VX_cluster.sv:88:5
				VX_pipe_register #(
					.DATAW(1),
					.RESETW(1),
					.DEPTH(1'd0)
				) __busy__(
					.clk(clk),
					.reset(reset),
					.enable(1'b1),
					.data_in(|per_socket_busy),
					.data_out(busy)
				);
			end
			assign cluster.clk = clk;
			assign cluster.reset = cluster_reset;
			assign per_cluster_busy[cluster_id] = cluster.busy;
		end
	endgenerate
	// Trace: src/Vortex.sv:117:5
	VX_pipe_register #(
		.DATAW(1),
		.RESETW(1),
		.DEPTH(1'd0)
	) __busy__(
		.clk(clk),
		.reset(reset),
		.enable(1'b1),
		.data_in(|per_cluster_busy),
		.data_out(busy)
	);
	// Trace: src/Vortex.sv:128:5
endmodule
// removed interface: VX_dispatch_if
module VX_mux (
	data_in,
	sel_in,
	data_out
);
	// Trace: src/VX_mux.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_mux.sv:3:15
	parameter N = 1;
	// Trace: src/VX_mux.sv:4:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_mux.sv:6:5
	input wire [(N * DATAW) - 1:0] data_in;
	// Trace: src/VX_mux.sv:7:5
	input wire [LN - 1:0] sel_in;
	// Trace: src/VX_mux.sv:8:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_mux.sv:10:5
	generate
		if (N > 1) begin : g_mux
			// Trace: src/VX_mux.sv:11:9
			assign data_out = data_in[sel_in * DATAW+:DATAW];
		end
		else begin : g_passthru
			// Trace: src/VX_mux.sv:13:9
			assign data_out = data_in;
		end
	endgenerate
endmodule
module VX_onehot_encoder (
	data_in,
	data_out,
	valid_out
);
	// Trace: src/VX_onehot_encoder.sv:2:15
	parameter N = 1;
	// Trace: src/VX_onehot_encoder.sv:3:15
	parameter REVERSE = 0;
	// Trace: src/VX_onehot_encoder.sv:4:15
	parameter MODEL = 1;
	// Trace: src/VX_onehot_encoder.sv:5:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_onehot_encoder.sv:7:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_onehot_encoder.sv:8:5
	output wire [LN - 1:0] data_out;
	// Trace: src/VX_onehot_encoder.sv:9:5
	output wire valid_out;
	// Trace: src/VX_onehot_encoder.sv:11:5
	function automatic signed [LN - 1:0] sv2v_cast_83428_signed;
		input reg signed [LN - 1:0] inp;
		sv2v_cast_83428_signed = inp;
	endfunction
	generate
		if (N == 1) begin : g_n1
			// Trace: src/VX_onehot_encoder.sv:12:9
			assign data_out = 0;
			// Trace: src/VX_onehot_encoder.sv:13:9
			assign valid_out = data_in;
		end
		else if (N == 2) begin : g_n2
			// Trace: src/VX_onehot_encoder.sv:15:9
			assign data_out = data_in[!REVERSE];
			// Trace: src/VX_onehot_encoder.sv:16:9
			assign valid_out = |data_in;
		end
		else if (MODEL == 1) begin : g_model1
			// Trace: src/VX_onehot_encoder.sv:18:9
			localparam M = 1 << LN;
			// Trace: src/VX_onehot_encoder.sv:19:9
			wire [M - 1:0] addr [0:LN - 1];
			// Trace: src/VX_onehot_encoder.sv:20:9
			wire [M - 1:0] v [0:LN + 0];
			// Trace: src/VX_onehot_encoder.sv:21:9
			function automatic [M - 1:0] sv2v_cast_ABEB2;
				input reg [M - 1:0] inp;
				sv2v_cast_ABEB2 = inp;
			endfunction
			assign v[0] = (REVERSE ? sv2v_cast_ABEB2(data_in) << (M - N) : sv2v_cast_ABEB2(data_in));
			genvar _gv_lvl_1;
			for (_gv_lvl_1 = 1; _gv_lvl_1 < (LN + 1); _gv_lvl_1 = _gv_lvl_1 + 1) begin : g_scan_l
				localparam lvl = _gv_lvl_1;
				// Trace: src/VX_onehot_encoder.sv:23:13
				localparam SN = 1 << (LN - lvl);
				// Trace: src/VX_onehot_encoder.sv:24:13
				localparam SI = M / SN;
				genvar _gv_s_1;
				for (_gv_s_1 = 0; _gv_s_1 < SN; _gv_s_1 = _gv_s_1 + 1) begin : g_scan_s
					localparam s = _gv_s_1;
					// Trace: src/VX_onehot_encoder.sv:26:17
					wire [1:0] vs = {v[lvl - 1][(s * SI) + (SI >> 1)], v[lvl - 1][s * SI]};
					// Trace: src/VX_onehot_encoder.sv:27:17
					assign v[lvl][s * SI] = |vs;
					if (lvl == 1) begin : g_lvl_1
						// Trace: src/VX_onehot_encoder.sv:29:21
						assign addr[lvl - 1][s * SI+:lvl] = vs[!REVERSE];
					end
					else begin : g_lvl_n
						// Trace: src/VX_onehot_encoder.sv:31:21
						assign addr[lvl - 1][s * SI+:lvl] = {vs[!REVERSE], addr[lvl - 2][s * SI+:lvl - 1] | addr[lvl - 2][(s * SI) + (SI >> 1)+:lvl - 1]};
					end
				end
			end
			// Trace: src/VX_onehot_encoder.sv:38:9
			assign data_out = addr[LN - 1][LN - 1:0];
			// Trace: src/VX_onehot_encoder.sv:39:9
			assign valid_out = v[LN][0];
		end
		else if ((MODEL == 2) && (REVERSE == 0)) begin : g_model2
			genvar _gv_j_16;
			for (_gv_j_16 = 0; _gv_j_16 < LN; _gv_j_16 = _gv_j_16 + 1) begin : g_data_out
				localparam j = _gv_j_16;
				// Trace: src/VX_onehot_encoder.sv:42:13
				wire [N - 1:0] mask;
				genvar _gv_i_134;
				for (_gv_i_134 = 0; _gv_i_134 < N; _gv_i_134 = _gv_i_134 + 1) begin : g_mask
					localparam i = _gv_i_134;
					// Trace: src/VX_onehot_encoder.sv:44:17
					assign mask[i] = i[j];
				end
				// Trace: src/VX_onehot_encoder.sv:46:13
				assign data_out[j] = |(mask & data_in);
			end
			// Trace: src/VX_onehot_encoder.sv:48:9
			assign valid_out = |data_in;
		end
		else begin : g_model0
			// Trace: src/VX_onehot_encoder.sv:50:9
			reg [LN - 1:0] index_w;
			if (REVERSE != 0) begin : g_msb
				// Trace: src/VX_onehot_encoder.sv:52:13
				always @(*) begin
					// Trace: src/VX_onehot_encoder.sv:53:17
					index_w = 1'sbx;
					// Trace: src/VX_onehot_encoder.sv:54:17
					begin : sv2v_autoblock_1
						// Trace: src/VX_onehot_encoder.sv:54:22
						integer i;
						// Trace: src/VX_onehot_encoder.sv:54:22
						for (i = N - 1; i >= 0; i = i - 1)
							begin
								// Trace: src/VX_onehot_encoder.sv:55:21
								if (data_in[i])
									// Trace: src/VX_onehot_encoder.sv:56:25
									index_w = sv2v_cast_83428_signed((N - 1) - i);
							end
					end
				end
			end
			else begin : g_lsb
				// Trace: src/VX_onehot_encoder.sv:61:13
				always @(*) begin
					// Trace: src/VX_onehot_encoder.sv:62:17
					index_w = 1'sbx;
					// Trace: src/VX_onehot_encoder.sv:63:17
					begin : sv2v_autoblock_2
						// Trace: src/VX_onehot_encoder.sv:63:22
						integer i;
						// Trace: src/VX_onehot_encoder.sv:63:22
						for (i = 0; i < N; i = i + 1)
							begin
								// Trace: src/VX_onehot_encoder.sv:64:21
								if (data_in[i])
									// Trace: src/VX_onehot_encoder.sv:65:25
									index_w = sv2v_cast_83428_signed(i);
							end
					end
				end
			end
			// Trace: src/VX_onehot_encoder.sv:70:9
			assign data_out = index_w;
			// Trace: src/VX_onehot_encoder.sv:71:9
			assign valid_out = |data_in;
		end
	endgenerate
endmodule
module VX_split_join (
	clk,
	reset,
	valid,
	wid,
	split,
	sjoin,
	join_valid,
	join_is_dvg,
	join_is_else,
	join_wid,
	join_tmask,
	join_pc,
	stack_wid,
	stack_ptr
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/VX_split_join.sv:2:16
	parameter INSTANCE_ID = "";
	// Trace: src/VX_split_join.sv:4:5
	input wire clk;
	// Trace: src/VX_split_join.sv:5:5
	input wire reset;
	// Trace: src/VX_split_join.sv:6:5
	input wire valid;
	// Trace: src/VX_split_join.sv:7:5
	input wire [1:0] wid;
	// Trace: src/VX_split_join.sv:8:5
	// removed localparam type VX_gpu_pkg_split_t
	input wire [40:0] split;
	// Trace: src/VX_split_join.sv:9:5
	// removed localparam type VX_gpu_pkg_join_t
	input wire [2:0] sjoin;
	// Trace: src/VX_split_join.sv:10:5
	output wire join_valid;
	// Trace: src/VX_split_join.sv:11:5
	output wire join_is_dvg;
	// Trace: src/VX_split_join.sv:12:5
	output wire join_is_else;
	// Trace: src/VX_split_join.sv:13:5
	output wire [1:0] join_wid;
	// Trace: src/VX_split_join.sv:14:5
	output wire [3:0] join_tmask;
	// Trace: src/VX_split_join.sv:15:5
	output wire [30:0] join_pc;
	// Trace: src/VX_split_join.sv:16:5
	input wire [1:0] stack_wid;
	// Trace: src/VX_split_join.sv:17:5
	output wire [1:0] stack_ptr;
	// Trace: src/VX_split_join.sv:19:5
	wire [34:0] ipdom_data [3:0];
	// Trace: src/VX_split_join.sv:20:5
	wire [1:0] ipdom_q_ptr [3:0];
	// Trace: src/VX_split_join.sv:21:5
	wire ipdom_set [3:0];
	// Trace: src/VX_split_join.sv:22:5
	wire [34:0] ipdom_q0 = {split[38-:4] | split[34-:4], 31'sd0};
	// Trace: src/VX_split_join.sv:23:5
	wire [34:0] ipdom_q1 = {split[34-:4], split[30-:31]};
	// Trace: src/VX_split_join.sv:24:5
	wire sjoin_is_dvg = sjoin[1-:2] != ipdom_q_ptr[wid];
	// Trace: src/VX_split_join.sv:25:5
	wire ipdom_push = (valid && split[40]) && split[39];
	// Trace: src/VX_split_join.sv:26:5
	wire ipdom_pop = (valid && sjoin[2]) && sjoin_is_dvg;
	// Trace: src/VX_split_join.sv:27:5
	genvar _gv_i_135;
	generate
		for (_gv_i_135 = 0; _gv_i_135 < 4; _gv_i_135 = _gv_i_135 + 1) begin : g_ipdom_stacks
			localparam i = _gv_i_135;
			// Trace: src/VX_split_join.sv:28:9
			VX_ipdom_stack #(
				.WIDTH(35),
				.DEPTH(3)
			) ipdom_stack(
				.clk(clk),
				.reset(reset),
				.q0(ipdom_q0),
				.q1(ipdom_q1),
				.d(ipdom_data[i]),
				.d_set(ipdom_set[i]),
				.q_ptr(ipdom_q_ptr[i]),
				.push(ipdom_push && (i == wid)),
				.pop(ipdom_pop && (i == wid)),
				.empty(),
				.full()
			);
		end
	endgenerate
	// Trace: src/VX_split_join.sv:45:5
	VX_pipe_register #(
		.DATAW(40),
		.DEPTH(1),
		.RESETW(1)
	) pipe_reg(
		.clk(clk),
		.reset(reset),
		.enable(1'b1),
		.data_in({valid && sjoin[2], sjoin_is_dvg, ipdom_set[wid], wid, ipdom_data[wid]}),
		.data_out({join_valid, join_is_dvg, join_is_else, join_wid, join_tmask, join_pc})
	);
	// Trace: src/VX_split_join.sv:56:5
	assign stack_ptr = ipdom_q_ptr[stack_wid];
endmodule
module VX_reduce (
	data_in,
	data_out
);
	// Trace: src/VX_reduce.sv:2:15
	parameter DATAW_IN = 1;
	// Trace: src/VX_reduce.sv:3:15
	parameter DATAW_OUT = DATAW_IN;
	// Trace: src/VX_reduce.sv:4:15
	parameter N = 1;
	// Trace: src/VX_reduce.sv:5:15
	parameter OP = "+";
	// Trace: src/VX_reduce.sv:7:5
	input wire [(N * DATAW_IN) - 1:0] data_in;
	// Trace: src/VX_reduce.sv:8:5
	output wire [DATAW_OUT - 1:0] data_out;
	// Trace: src/VX_reduce.sv:10:5
	function automatic [DATAW_OUT - 1:0] sv2v_cast_0EBAF;
		input reg [DATAW_OUT - 1:0] inp;
		sv2v_cast_0EBAF = inp;
	endfunction
	generate
		if (N == 1) begin : g_passthru
			// Trace: src/VX_reduce.sv:11:9
			assign data_out = sv2v_cast_0EBAF(data_in[0+:DATAW_IN]);
		end
		else begin : g_reduce
			// Trace: src/VX_reduce.sv:13:9
			localparam signed [31:0] N_A = N / 2;
			// Trace: src/VX_reduce.sv:14:9
			localparam signed [31:0] N_B = N - N_A;
			// Trace: src/VX_reduce.sv:15:9
			wire [(N_A * DATAW_IN) - 1:0] in_A;
			// Trace: src/VX_reduce.sv:16:9
			wire [(N_B * DATAW_IN) - 1:0] in_B;
			// Trace: src/VX_reduce.sv:17:9
			wire [DATAW_OUT - 1:0] out_A;
			wire [DATAW_OUT - 1:0] out_B;
			genvar _gv_i_136;
			for (_gv_i_136 = 0; _gv_i_136 < N_A; _gv_i_136 = _gv_i_136 + 1) begin : g_in_A
				localparam i = _gv_i_136;
				// Trace: src/VX_reduce.sv:19:13
				assign in_A[i * DATAW_IN+:DATAW_IN] = data_in[i * DATAW_IN+:DATAW_IN];
			end
			genvar _gv_i_137;
			for (_gv_i_137 = 0; _gv_i_137 < N_B; _gv_i_137 = _gv_i_137 + 1) begin : g_in_B
				localparam i = _gv_i_137;
				// Trace: src/VX_reduce.sv:22:13
				assign in_B[i * DATAW_IN+:DATAW_IN] = data_in[(N_A + i) * DATAW_IN+:DATAW_IN];
			end
			// Trace: src/VX_reduce.sv:24:9
			VX_reduce #(
				.DATAW_IN(DATAW_IN),
				.DATAW_OUT(DATAW_OUT),
				.N(N_A),
				.OP(OP)
			) reduce_A(
				.data_in(in_A),
				.data_out(out_A)
			);
			// Trace: src/VX_reduce.sv:33:9
			VX_reduce #(
				.DATAW_IN(DATAW_IN),
				.DATAW_OUT(DATAW_OUT),
				.N(N_B),
				.OP(OP)
			) reduce_B(
				.data_in(in_B),
				.data_out(out_B)
			);
			if (OP == "+") begin : g_plus
				// Trace: src/VX_reduce.sv:43:13
				assign data_out = out_A + out_B;
			end
			else if (OP == "^") begin : g_xor
				// Trace: src/VX_reduce.sv:45:13
				assign data_out = out_A ^ out_B;
			end
			else if (OP == "&") begin : g_and
				// Trace: src/VX_reduce.sv:47:13
				assign data_out = out_A & out_B;
			end
			else if (OP == "|") begin : g_or
				// Trace: src/VX_reduce.sv:49:13
				assign data_out = out_A | out_B;
			end
		end
	endgenerate
endmodule
module VX_scan (
	data_in,
	data_out
);
	// Trace: src/VX_scan.sv:2:15
	parameter N = 1;
	// Trace: src/VX_scan.sv:3:15
	parameter OP = "^";
	// Trace: src/VX_scan.sv:4:15
	parameter REVERSE = 0;
	// Trace: src/VX_scan.sv:6:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_scan.sv:7:5
	output wire [N - 1:0] data_out;
	// Trace: src/VX_scan.sv:9:5
	localparam LOGN = $clog2(N);
	// Trace: src/VX_scan.sv:10:5
	wire [(LOGN >= 0 ? ((LOGN + 1) * N) - 1 : ((1 - LOGN) * N) + ((LOGN * N) - 1)):(LOGN >= 0 ? 0 : LOGN * N)] t;
	// Trace: src/VX_scan.sv:11:5
	generate
		if (REVERSE != 0) begin : g_data_in_reverse
			// Trace: src/VX_scan.sv:12:9
			assign t[(LOGN >= 0 ? 0 : LOGN) * N+:N] = data_in;
		end
		else begin : g_data_in_no_reverse
			// Trace: src/VX_scan.sv:14:9
			function automatic [N - 1:0] _sv2v_strm_F2A76;
				input reg [(0 + N) - 1:0] inp;
				reg [(0 + N) - 1:0] _sv2v_strm_55E18_inp;
				reg [(0 + N) - 1:0] _sv2v_strm_55E18_out;
				integer _sv2v_strm_55E18_idx;
				begin
					_sv2v_strm_55E18_inp = {inp};
					for (_sv2v_strm_55E18_idx = 0; _sv2v_strm_55E18_idx <= ((0 + N) - 1); _sv2v_strm_55E18_idx = _sv2v_strm_55E18_idx + 1)
						_sv2v_strm_55E18_out[((0 + N) - 1) - _sv2v_strm_55E18_idx-:1] = _sv2v_strm_55E18_inp[_sv2v_strm_55E18_idx+:1];
					_sv2v_strm_F2A76 = ((0 + N) <= N ? _sv2v_strm_55E18_out << (N - (0 + N)) : _sv2v_strm_55E18_out >> ((0 + N) - N));
				end
			endfunction
			assign t[(LOGN >= 0 ? 0 : LOGN) * N+:N] = _sv2v_strm_F2A76({data_in});
		end
	endgenerate
	// Trace: src/VX_scan.sv:16:5
	function automatic [N - 1:0] sv2v_cast_AC047;
		input reg [N - 1:0] inp;
		sv2v_cast_AC047 = inp;
	endfunction
	generate
		if ((N == 2) && (OP == "&")) begin : g_scan_n2_and
			// Trace: src/VX_scan.sv:17:6
			assign t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N] = {t[((LOGN >= 0 ? 0 : LOGN) * N) + 1], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 1-:2]};
		end
		else if ((N == 3) && (OP == "&")) begin : g_scan_n3_and
			// Trace: src/VX_scan.sv:19:6
			assign t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N] = {t[((LOGN >= 0 ? 0 : LOGN) * N) + 2], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 2-:2], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 2-:3]};
		end
		else if ((N == 4) && (OP == "&")) begin : g_scan_n4_and
			// Trace: src/VX_scan.sv:21:6
			assign t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N] = {t[((LOGN >= 0 ? 0 : LOGN) * N) + 3], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 3-:2], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 3-:3], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 3-:4]};
		end
		else begin : g_scan
			// Trace: src/VX_scan.sv:23:9
			wire [N - 1:0] fill;
			genvar _gv_i_138;
			for (_gv_i_138 = 0; _gv_i_138 < LOGN; _gv_i_138 = _gv_i_138 + 1) begin : g_i
				localparam i = _gv_i_138;
				// Trace: src/VX_scan.sv:25:13
				wire [N - 1:0] shifted = sv2v_cast_AC047({fill, t[(LOGN >= 0 ? i : LOGN - i) * N+:N]} >> (1 << i));
				if (OP == "^") begin : g_xor
					// Trace: src/VX_scan.sv:27:11
					assign fill = {N {1'b0}};
					// Trace: src/VX_scan.sv:28:11
					assign t[(LOGN >= 0 ? i + 1 : LOGN - (i + 1)) * N+:N] = t[(LOGN >= 0 ? i : LOGN - i) * N+:N] ^ shifted;
				end
				else if (OP == "&") begin : g_and
					// Trace: src/VX_scan.sv:30:11
					assign fill = {N {1'b1}};
					// Trace: src/VX_scan.sv:31:11
					assign t[(LOGN >= 0 ? i + 1 : LOGN - (i + 1)) * N+:N] = t[(LOGN >= 0 ? i : LOGN - i) * N+:N] & shifted;
				end
				else if (OP == "|") begin : g_or
					// Trace: src/VX_scan.sv:33:11
					assign fill = {N {1'b0}};
					// Trace: src/VX_scan.sv:34:11
					assign t[(LOGN >= 0 ? i + 1 : LOGN - (i + 1)) * N+:N] = t[(LOGN >= 0 ? i : LOGN - i) * N+:N] | shifted;
				end
			end
		end
	endgenerate
	// Trace: src/VX_scan.sv:38:5
	generate
		if (REVERSE != 0) begin : g_data_out_reverse
			// Trace: src/VX_scan.sv:39:9
			assign data_out = t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N];
		end
		else begin : g_data_out
			genvar _gv_i_139;
			for (_gv_i_139 = 0; _gv_i_139 < N; _gv_i_139 = _gv_i_139 + 1) begin : g_i
				localparam i = _gv_i_139;
				// Trace: src/VX_scan.sv:42:13
				assign data_out[i] = t[((LOGN >= 0 ? LOGN : LOGN - LOGN) * N) + ((N - 1) - i)];
			end
		end
	endgenerate
endmodule
module VX_priority_encoder (
	data_in,
	onehot_out,
	index_out,
	valid_out
);
	// Trace: src/VX_priority_encoder.sv:2:15
	parameter N = 1;
	// Trace: src/VX_priority_encoder.sv:3:15
	parameter REVERSE = 0;
	// Trace: src/VX_priority_encoder.sv:4:15
	parameter MODEL = 1;
	// Trace: src/VX_priority_encoder.sv:5:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_priority_encoder.sv:7:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_priority_encoder.sv:8:5
	output wire [N - 1:0] onehot_out;
	// Trace: src/VX_priority_encoder.sv:9:5
	output wire [LN - 1:0] index_out;
	// Trace: src/VX_priority_encoder.sv:10:5
	output wire valid_out;
	// Trace: src/VX_priority_encoder.sv:12:5
	wire [N - 1:0] reversed;
	// Trace: src/VX_priority_encoder.sv:13:5
	generate
		if (REVERSE != 0) begin : g_reverse
			genvar _gv_i_140;
			for (_gv_i_140 = 0; _gv_i_140 < N; _gv_i_140 = _gv_i_140 + 1) begin : g_i
				localparam i = _gv_i_140;
				// Trace: src/VX_priority_encoder.sv:15:13
				assign reversed[(N - i) - 1] = data_in[i];
			end
		end
		else begin : g_no_reverse
			// Trace: src/VX_priority_encoder.sv:18:9
			assign reversed = data_in;
		end
	endgenerate
	// Trace: src/VX_priority_encoder.sv:20:5
	function automatic signed [LN - 1:0] sv2v_cast_83428_signed;
		input reg signed [LN - 1:0] inp;
		sv2v_cast_83428_signed = inp;
	endfunction
	function automatic signed [N - 1:0] sv2v_cast_AC047_signed;
		input reg signed [N - 1:0] inp;
		sv2v_cast_AC047_signed = inp;
	endfunction
	generate
		if (N == 1) begin : g_n1
			// Trace: src/VX_priority_encoder.sv:21:9
			assign onehot_out = reversed;
			// Trace: src/VX_priority_encoder.sv:22:9
			assign index_out = 1'sb0;
			// Trace: src/VX_priority_encoder.sv:23:9
			assign valid_out = reversed;
		end
		else if (N == 2) begin : g_n2
			// Trace: src/VX_priority_encoder.sv:25:9
			assign onehot_out = {reversed[1] && ~reversed[0], reversed[0]};
			// Trace: src/VX_priority_encoder.sv:26:9
			assign index_out = ~reversed[0];
			// Trace: src/VX_priority_encoder.sv:27:9
			assign valid_out = |reversed;
		end
		else if (MODEL == 1) begin : g_model1
			// Trace: src/VX_priority_encoder.sv:29:9
			wire [N - 1:0] higher_pri_regs;
			// Trace: src/VX_priority_encoder.sv:30:9
			assign higher_pri_regs[0] = 1'b0;
			genvar _gv_i_141;
			for (_gv_i_141 = 1; _gv_i_141 < N; _gv_i_141 = _gv_i_141 + 1) begin : g_higher_pri_regs
				localparam i = _gv_i_141;
				// Trace: src/VX_priority_encoder.sv:32:13
				assign higher_pri_regs[i] = higher_pri_regs[i - 1] | reversed[i - 1];
			end
			// Trace: src/VX_priority_encoder.sv:34:9
			assign onehot_out[N - 1:0] = reversed[N - 1:0] & ~higher_pri_regs[N - 1:0];
			// Trace: src/VX_priority_encoder.sv:35:9
			VX_lzc #(
				.N(N),
				.REVERSE(1)
			) lzc(
				.data_in(reversed),
				.data_out(index_out),
				.valid_out(valid_out)
			);
		end
		else if (MODEL == 2) begin : g_model2
			// Trace: src/VX_priority_encoder.sv:44:9
			wire [N - 1:0] scan_lo;
			// Trace: src/VX_priority_encoder.sv:45:9
			VX_scan #(
				.N(N),
				.OP("|")
			) scan(
				.data_in(reversed),
				.data_out(scan_lo)
			);
			// Trace: src/VX_priority_encoder.sv:52:9
			VX_lzc #(
				.N(N),
				.REVERSE(1)
			) lzc(
				.data_in(reversed),
				.data_out(index_out),
				.valid_out(valid_out)
			);
			// Trace: src/VX_priority_encoder.sv:60:9
			assign onehot_out = scan_lo & {~scan_lo[N - 2:0], 1'b1};
		end
		else if (MODEL == 3) begin : g_model3
			// Trace: src/VX_priority_encoder.sv:62:9
			assign onehot_out = reversed & -reversed;
			// Trace: src/VX_priority_encoder.sv:63:9
			VX_lzc #(
				.N(N),
				.REVERSE(1)
			) lzc(
				.data_in(reversed),
				.data_out(index_out),
				.valid_out(valid_out)
			);
		end
		else begin : g_model0
			// Trace: src/VX_priority_encoder.sv:72:9
			reg [LN - 1:0] index_w;
			// Trace: src/VX_priority_encoder.sv:73:9
			reg [N - 1:0] onehot_w;
			// Trace: src/VX_priority_encoder.sv:74:9
			always @(*) begin
				// Trace: src/VX_priority_encoder.sv:75:13
				index_w = 1'sbx;
				// Trace: src/VX_priority_encoder.sv:76:13
				onehot_w = 1'sbx;
				// Trace: src/VX_priority_encoder.sv:77:13
				begin : sv2v_autoblock_1
					// Trace: src/VX_priority_encoder.sv:77:18
					integer i;
					// Trace: src/VX_priority_encoder.sv:77:18
					for (i = N - 1; i >= 0; i = i - 1)
						begin
							// Trace: src/VX_priority_encoder.sv:78:17
							if (reversed[i]) begin
								// Trace: src/VX_priority_encoder.sv:79:21
								index_w = sv2v_cast_83428_signed(i);
								// Trace: src/VX_priority_encoder.sv:80:21
								onehot_w = sv2v_cast_AC047_signed(1) << i;
							end
						end
				end
			end
			// Trace: src/VX_priority_encoder.sv:84:9
			assign index_out = index_w;
			// Trace: src/VX_priority_encoder.sv:85:9
			assign onehot_out = onehot_w;
			// Trace: src/VX_priority_encoder.sv:86:9
			assign valid_out = |reversed;
		end
	endgenerate
endmodule
module VX_reset_relay (
	clk,
	reset,
	reset_o
);
	// Trace: src/VX_reset_relay.sv:2:15
	parameter N = 1;
	// Trace: src/VX_reset_relay.sv:3:15
	parameter MAX_FANOUT = 0;
	// Trace: src/VX_reset_relay.sv:5:5
	input wire clk;
	// Trace: src/VX_reset_relay.sv:6:5
	input wire reset;
	// Trace: src/VX_reset_relay.sv:7:5
	output wire [N - 1:0] reset_o;
	// Trace: src/VX_reset_relay.sv:9:5
	generate
		if ((MAX_FANOUT >= 0) && (N > (MAX_FANOUT + (MAX_FANOUT / 2)))) begin : g_relay
			// Trace: src/VX_reset_relay.sv:10:9
			localparam F = (MAX_FANOUT > 0 ? MAX_FANOUT : 1);
			// Trace: src/VX_reset_relay.sv:11:9
			localparam R = N / F;
			// Trace: src/VX_reset_relay.sv:12:10
			reg [R - 1:0] reset_r;
			genvar _gv_i_142;
			for (_gv_i_142 = 0; _gv_i_142 < R; _gv_i_142 = _gv_i_142 + 1) begin : g_reset_r
				localparam i = _gv_i_142;
				// Trace: src/VX_reset_relay.sv:14:13
				always @(posedge clk)
					// Trace: src/VX_reset_relay.sv:15:17
					reset_r[i] <= reset;
			end
			genvar _gv_i_143;
			for (_gv_i_143 = 0; _gv_i_143 < N; _gv_i_143 = _gv_i_143 + 1) begin : g_reset_o
				localparam i = _gv_i_143;
				// Trace: src/VX_reset_relay.sv:19:13
				assign reset_o[i] = reset_r[i / F];
			end
		end
		else begin : g_passthru
			// Trace: src/VX_reset_relay.sv:22:9
			assign reset_o = {N {reset}};
		end
	endgenerate
endmodule
module VX_cache_mshr (
	clk,
	reset,
	deq_req_uuid,
	alc_req_uuid,
	fin_req_uuid,
	fill_valid,
	fill_id,
	fill_addr,
	dequeue_valid,
	dequeue_addr,
	dequeue_rw,
	dequeue_data,
	dequeue_id,
	dequeue_ready,
	allocate_valid,
	allocate_addr,
	allocate_rw,
	allocate_data,
	allocate_id,
	allocate_pending,
	allocate_previd,
	allocate_ready,
	finalize_valid,
	finalize_is_release,
	finalize_is_pending,
	finalize_previd,
	finalize_id
);
	// Trace: src/VX_cache_mshr.sv:2:16
	parameter INSTANCE_ID = "";
	// Trace: src/VX_cache_mshr.sv:3:15
	parameter BANK_ID = 0;
	// Trace: src/VX_cache_mshr.sv:4:15
	parameter LINE_SIZE = 16;
	// Trace: src/VX_cache_mshr.sv:5:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_mshr.sv:6:15
	parameter MSHR_SIZE = 4;
	// Trace: src/VX_cache_mshr.sv:7:15
	parameter UUID_WIDTH = 0;
	// Trace: src/VX_cache_mshr.sv:8:15
	parameter DATA_WIDTH = 1;
	// Trace: src/VX_cache_mshr.sv:9:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_cache_mshr.sv:10:15
	parameter MSHR_ADDR_WIDTH = (MSHR_SIZE > 1 ? $clog2(MSHR_SIZE) : 1);
	// Trace: src/VX_cache_mshr.sv:12:5
	input wire clk;
	// Trace: src/VX_cache_mshr.sv:13:5
	input wire reset;
	// Trace: src/VX_cache_mshr.sv:14:5
	input wire [(UUID_WIDTH > 0 ? UUID_WIDTH : 1) - 1:0] deq_req_uuid;
	// Trace: src/VX_cache_mshr.sv:15:5
	input wire [(UUID_WIDTH > 0 ? UUID_WIDTH : 1) - 1:0] alc_req_uuid;
	// Trace: src/VX_cache_mshr.sv:16:5
	input wire [(UUID_WIDTH > 0 ? UUID_WIDTH : 1) - 1:0] fin_req_uuid;
	// Trace: src/VX_cache_mshr.sv:17:5
	input wire fill_valid;
	// Trace: src/VX_cache_mshr.sv:18:5
	input wire [MSHR_ADDR_WIDTH - 1:0] fill_id;
	// Trace: src/VX_cache_mshr.sv:19:5
	output wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] fill_addr;
	// Trace: src/VX_cache_mshr.sv:20:5
	output wire dequeue_valid;
	// Trace: src/VX_cache_mshr.sv:21:5
	output wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] dequeue_addr;
	// Trace: src/VX_cache_mshr.sv:22:5
	output wire dequeue_rw;
	// Trace: src/VX_cache_mshr.sv:23:5
	output wire [DATA_WIDTH - 1:0] dequeue_data;
	// Trace: src/VX_cache_mshr.sv:24:5
	output wire [MSHR_ADDR_WIDTH - 1:0] dequeue_id;
	// Trace: src/VX_cache_mshr.sv:25:5
	input wire dequeue_ready;
	// Trace: src/VX_cache_mshr.sv:26:5
	input wire allocate_valid;
	// Trace: src/VX_cache_mshr.sv:27:5
	input wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] allocate_addr;
	// Trace: src/VX_cache_mshr.sv:28:5
	input wire allocate_rw;
	// Trace: src/VX_cache_mshr.sv:29:5
	input wire [DATA_WIDTH - 1:0] allocate_data;
	// Trace: src/VX_cache_mshr.sv:30:5
	output wire [MSHR_ADDR_WIDTH - 1:0] allocate_id;
	// Trace: src/VX_cache_mshr.sv:31:5
	output wire allocate_pending;
	// Trace: src/VX_cache_mshr.sv:32:5
	output wire [MSHR_ADDR_WIDTH - 1:0] allocate_previd;
	// Trace: src/VX_cache_mshr.sv:33:5
	output wire allocate_ready;
	// Trace: src/VX_cache_mshr.sv:34:5
	input wire finalize_valid;
	// Trace: src/VX_cache_mshr.sv:35:5
	input wire finalize_is_release;
	// Trace: src/VX_cache_mshr.sv:36:5
	input wire finalize_is_pending;
	// Trace: src/VX_cache_mshr.sv:37:5
	input wire [MSHR_ADDR_WIDTH - 1:0] finalize_previd;
	// Trace: src/VX_cache_mshr.sv:38:5
	input wire [MSHR_ADDR_WIDTH - 1:0] finalize_id;
	// Trace: src/VX_cache_mshr.sv:40:5
	reg [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_table [0:MSHR_SIZE - 1];
	// Trace: src/VX_cache_mshr.sv:41:5
	reg [MSHR_ADDR_WIDTH - 1:0] next_index [0:MSHR_SIZE - 1];
	// Trace: src/VX_cache_mshr.sv:42:5
	reg [MSHR_SIZE - 1:0] valid_table;
	reg [MSHR_SIZE - 1:0] valid_table_n;
	// Trace: src/VX_cache_mshr.sv:43:5
	reg [MSHR_SIZE - 1:0] next_table;
	reg [MSHR_SIZE - 1:0] next_table_x;
	reg [MSHR_SIZE - 1:0] next_table_n;
	// Trace: src/VX_cache_mshr.sv:44:5
	reg [MSHR_SIZE - 1:0] write_table;
	// Trace: src/VX_cache_mshr.sv:45:5
	reg allocate_rdy;
	reg allocate_rdy_n;
	// Trace: src/VX_cache_mshr.sv:46:5
	reg [MSHR_ADDR_WIDTH - 1:0] allocate_id_r;
	reg [MSHR_ADDR_WIDTH - 1:0] allocate_id_n;
	// Trace: src/VX_cache_mshr.sv:47:5
	reg dequeue_val;
	reg dequeue_val_n;
	// Trace: src/VX_cache_mshr.sv:48:5
	reg [MSHR_ADDR_WIDTH - 1:0] dequeue_id_r;
	reg [MSHR_ADDR_WIDTH - 1:0] dequeue_id_n;
	// Trace: src/VX_cache_mshr.sv:49:5
	wire [MSHR_ADDR_WIDTH - 1:0] prev_idx;
	// Trace: src/VX_cache_mshr.sv:50:5
	wire allocate_fire = allocate_valid && allocate_ready;
	// Trace: src/VX_cache_mshr.sv:51:5
	wire dequeue_fire = dequeue_valid && dequeue_ready;
	// Trace: src/VX_cache_mshr.sv:52:5
	wire [MSHR_SIZE - 1:0] addr_matches;
	// Trace: src/VX_cache_mshr.sv:53:5
	genvar _gv_i_144;
	generate
		for (_gv_i_144 = 0; _gv_i_144 < MSHR_SIZE; _gv_i_144 = _gv_i_144 + 1) begin : g_addr_matches
			localparam i = _gv_i_144;
			// Trace: src/VX_cache_mshr.sv:54:9
			assign addr_matches[i] = valid_table[i] && (addr_table[i] == allocate_addr);
		end
	endgenerate
	// Trace: src/VX_cache_mshr.sv:56:5
	// rewrote reg-to-output bindings
	wire [MSHR_ADDR_WIDTH:1] sv2v_tmp_allocate_sel_data_out;
	always @(*) allocate_id_n = sv2v_tmp_allocate_sel_data_out;
	wire [1:1] sv2v_tmp_allocate_sel_valid_out;
	always @(*) allocate_rdy_n = sv2v_tmp_allocate_sel_valid_out;
	VX_lzc #(
		.N(MSHR_SIZE),
		.REVERSE(1)
	) allocate_sel(
		.data_in(~valid_table_n),
		.data_out(sv2v_tmp_allocate_sel_data_out),
		.valid_out(sv2v_tmp_allocate_sel_valid_out)
	);
	// Trace: src/VX_cache_mshr.sv:64:5
	VX_priority_encoder #(.N(MSHR_SIZE)) prev_sel(
		.data_in(addr_matches & ~next_table_x),
		.index_out(prev_idx),
		.onehot_out(),
		.valid_out()
	);
	// Trace: src/VX_cache_mshr.sv:72:5
	always @(*) begin
		// Trace: src/VX_cache_mshr.sv:73:9
		valid_table_n = valid_table;
		// Trace: src/VX_cache_mshr.sv:74:9
		next_table_x = next_table;
		// Trace: src/VX_cache_mshr.sv:75:9
		dequeue_val_n = dequeue_val;
		// Trace: src/VX_cache_mshr.sv:76:9
		dequeue_id_n = dequeue_id;
		// Trace: src/VX_cache_mshr.sv:77:9
		if (fill_valid) begin
			// Trace: src/VX_cache_mshr.sv:78:13
			dequeue_val_n = 1;
			// Trace: src/VX_cache_mshr.sv:79:13
			dequeue_id_n = fill_id;
		end
		if (dequeue_fire) begin
			// Trace: src/VX_cache_mshr.sv:82:13
			valid_table_n[dequeue_id] = 0;
			// Trace: src/VX_cache_mshr.sv:83:13
			if (next_table[dequeue_id])
				// Trace: src/VX_cache_mshr.sv:84:17
				dequeue_id_n = next_index[dequeue_id];
			else if ((finalize_valid && finalize_is_pending) && (finalize_previd == dequeue_id))
				// Trace: src/VX_cache_mshr.sv:86:17
				dequeue_id_n = finalize_id;
			else
				// Trace: src/VX_cache_mshr.sv:88:17
				dequeue_val_n = 0;
		end
		if (finalize_valid) begin
			// Trace: src/VX_cache_mshr.sv:92:13
			if (finalize_is_release)
				// Trace: src/VX_cache_mshr.sv:93:17
				valid_table_n[finalize_id] = 0;
			if (finalize_is_pending)
				// Trace: src/VX_cache_mshr.sv:96:17
				next_table_x[finalize_previd] = 1;
		end
		// Trace: src/VX_cache_mshr.sv:99:9
		next_table_n = next_table_x;
		if (allocate_fire) begin
			// Trace: src/VX_cache_mshr.sv:101:13
			valid_table_n[allocate_id] = 1;
			// Trace: src/VX_cache_mshr.sv:102:13
			next_table_n[allocate_id] = 0;
		end
	end
	// Trace: src/VX_cache_mshr.sv:105:5
	always @(posedge clk) begin
		// Trace: src/VX_cache_mshr.sv:106:9
		if (reset) begin
			// Trace: src/VX_cache_mshr.sv:107:13
			valid_table <= 1'sb0;
			// Trace: src/VX_cache_mshr.sv:108:13
			allocate_rdy <= 0;
			// Trace: src/VX_cache_mshr.sv:109:13
			dequeue_val <= 0;
		end
		else begin
			// Trace: src/VX_cache_mshr.sv:111:13
			valid_table <= valid_table_n;
			// Trace: src/VX_cache_mshr.sv:112:13
			allocate_rdy <= allocate_rdy_n;
			// Trace: src/VX_cache_mshr.sv:113:13
			dequeue_val <= dequeue_val_n;
		end
		if (allocate_fire) begin
			// Trace: src/VX_cache_mshr.sv:116:13
			addr_table[allocate_id] <= allocate_addr;
			// Trace: src/VX_cache_mshr.sv:117:13
			write_table[allocate_id] <= allocate_rw;
		end
		if (finalize_valid && finalize_is_pending)
			// Trace: src/VX_cache_mshr.sv:120:13
			next_index[finalize_previd] <= finalize_id;
		// Trace: src/VX_cache_mshr.sv:122:9
		dequeue_id_r <= dequeue_id_n;
		// Trace: src/VX_cache_mshr.sv:123:9
		allocate_id_r <= allocate_id_n;
		// Trace: src/VX_cache_mshr.sv:124:9
		next_table <= next_table_n;
	end
	// Trace: src/VX_cache_mshr.sv:126:5
	VX_dp_ram #(
		.DATAW(DATA_WIDTH),
		.SIZE(MSHR_SIZE),
		.RDW_MODE("R"),
		.RADDR_REG(1)
	) mshr_store(
		.clk(clk),
		.reset(reset),
		.read(1'b1),
		.write(allocate_valid),
		.wren(1'b1),
		.waddr(allocate_id_r),
		.wdata(allocate_data),
		.raddr(dequeue_id_r),
		.rdata(dequeue_data)
	);
	// Trace: src/VX_cache_mshr.sv:142:5
	assign fill_addr = addr_table[fill_id];
	// Trace: src/VX_cache_mshr.sv:143:5
	assign allocate_ready = allocate_rdy;
	// Trace: src/VX_cache_mshr.sv:144:5
	assign allocate_id = allocate_id_r;
	// Trace: src/VX_cache_mshr.sv:145:5
	assign allocate_previd = prev_idx;
	// Trace: src/VX_cache_mshr.sv:146:5
	generate
		if (WRITEBACK) begin : g_pending_wb
			// Trace: src/VX_cache_mshr.sv:147:9
			assign allocate_pending = |addr_matches;
		end
		else begin : g_pending_wt
			// Trace: src/VX_cache_mshr.sv:149:9
			assign allocate_pending = |(addr_matches & ~write_table);
		end
	endgenerate
	// Trace: src/VX_cache_mshr.sv:151:5
	assign dequeue_valid = dequeue_val;
	// Trace: src/VX_cache_mshr.sv:152:5
	assign dequeue_addr = addr_table[dequeue_id_r];
	// Trace: src/VX_cache_mshr.sv:153:5
	assign dequeue_rw = write_table[dequeue_id_r];
	// Trace: src/VX_cache_mshr.sv:154:5
	assign dequeue_id = dequeue_id_r;
endmodule
// removed module with interface ports: VX_schedule
module VX_cyclic_arbiter (
	clk,
	reset,
	requests,
	grant_index,
	grant_onehot,
	grant_valid,
	grant_ready
);
	// Trace: src/VX_cyclic_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_cyclic_arbiter.sv:3:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_cyclic_arbiter.sv:5:5
	input wire clk;
	// Trace: src/VX_cyclic_arbiter.sv:6:5
	input wire reset;
	// Trace: src/VX_cyclic_arbiter.sv:7:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_cyclic_arbiter.sv:8:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_cyclic_arbiter.sv:9:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_cyclic_arbiter.sv:10:5
	output wire grant_valid;
	// Trace: src/VX_cyclic_arbiter.sv:11:5
	input wire grant_ready;
	// Trace: src/VX_cyclic_arbiter.sv:13:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_REQS == 1) begin : g_passthru
			// Trace: src/VX_cyclic_arbiter.sv:14:9
			assign grant_index = 1'sb0;
			// Trace: src/VX_cyclic_arbiter.sv:15:9
			assign grant_onehot = requests;
			// Trace: src/VX_cyclic_arbiter.sv:16:9
			assign grant_valid = requests[0];
		end
		else begin : g_arbiter
			// Trace: src/VX_cyclic_arbiter.sv:18:9
			localparam IS_POW2 = (1 << LOG_NUM_REQS) == NUM_REQS;
			// Trace: src/VX_cyclic_arbiter.sv:19:9
			wire [LOG_NUM_REQS - 1:0] grant_index_um;
			// Trace: src/VX_cyclic_arbiter.sv:20:9
			wire [NUM_REQS - 1:0] grant_onehot_w;
			wire [NUM_REQS - 1:0] grant_onehot_um;
			// Trace: src/VX_cyclic_arbiter.sv:21:9
			reg [LOG_NUM_REQS - 1:0] grant_index_r;
			// Trace: src/VX_cyclic_arbiter.sv:22:9
			always @(posedge clk)
				// Trace: src/VX_cyclic_arbiter.sv:23:13
				if (reset)
					// Trace: src/VX_cyclic_arbiter.sv:24:17
					grant_index_r <= 1'sb0;
				else if (grant_valid && grant_ready) begin
					begin
						// Trace: src/VX_cyclic_arbiter.sv:26:17
						if (!IS_POW2 && (grant_index == sv2v_cast_76B5F_signed(NUM_REQS - 1)))
							// Trace: src/VX_cyclic_arbiter.sv:27:21
							grant_index_r <= 1'sb0;
						else
							// Trace: src/VX_cyclic_arbiter.sv:29:21
							grant_index_r <= grant_index + sv2v_cast_76B5F_signed(1);
					end
				end
			// Trace: src/VX_cyclic_arbiter.sv:33:9
			VX_priority_encoder #(.N(NUM_REQS)) priority_encoder(
				.data_in(requests),
				.onehot_out(grant_onehot_um),
				.index_out(grant_index_um),
				.valid_out(grant_valid)
			);
			// Trace: src/VX_cyclic_arbiter.sv:41:9
			VX_demux #(
				.DATAW(1),
				.N(NUM_REQS)
			) grant_decoder(
				.sel_in(grant_index),
				.data_in(1'b1),
				.data_out(grant_onehot_w)
			);
			// Trace: src/VX_cyclic_arbiter.sv:49:9
			wire is_hit = requests[grant_index_r];
			// Trace: src/VX_cyclic_arbiter.sv:50:9
			assign grant_index = (is_hit ? grant_index_r : grant_index_um);
			// Trace: src/VX_cyclic_arbiter.sv:51:9
			assign grant_onehot = (is_hit ? grant_onehot_w : grant_onehot_um);
		end
	endgenerate
endmodule
module VX_demux (
	sel_in,
	data_in,
	data_out
);
	// Trace: src/VX_demux.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_demux.sv:3:15
	parameter N = 0;
	// Trace: src/VX_demux.sv:4:15
	parameter MODEL = 0;
	// Trace: src/VX_demux.sv:5:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_demux.sv:7:5
	input wire [LN - 1:0] sel_in;
	// Trace: src/VX_demux.sv:8:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_demux.sv:9:5
	output wire [(N * DATAW) - 1:0] data_out;
	// Trace: src/VX_demux.sv:11:5
	function automatic [(N * DATAW) - 1:0] sv2v_cast_3AE7C;
		input reg [(N * DATAW) - 1:0] inp;
		sv2v_cast_3AE7C = inp;
	endfunction
	generate
		if (N > 1) begin : g_demux
			// Trace: src/VX_demux.sv:12:9
			reg [(N * DATAW) - 1:0] shift;
			if (MODEL == 1) begin : g_model1
				// Trace: src/VX_demux.sv:14:13
				always @(*) begin
					// Trace: src/VX_demux.sv:15:17
					shift = 1'sb0;
					// Trace: src/VX_demux.sv:16:17
					shift[sel_in * DATAW+:DATAW] = {DATAW {1'b1}};
				end
			end
			else begin : g_model0
				// Trace: src/VX_demux.sv:19:13
				wire [N * DATAW:1] sv2v_tmp_6BA10;
				assign sv2v_tmp_6BA10 = sv2v_cast_3AE7C({DATAW {1'b1}}) << (sel_in * DATAW);
				always @(*) shift = sv2v_tmp_6BA10;
			end
			// Trace: src/VX_demux.sv:21:9
			assign data_out = {N {data_in}} & shift;
		end
		else begin : g_passthru
			// Trace: src/VX_demux.sv:23:9
			assign data_out = data_in;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_lsu_adapter
// removed module with interface ports: VX_dcr_data
// removed module with interface ports: VX_dispatch
// removed module with interface ports: VX_socket
// removed module with interface ports: VX_mem_switch
module VX_elastic_buffer (
	clk,
	reset,
	valid_in,
	ready_in,
	data_in,
	data_out,
	ready_out,
	valid_out
);
	// Trace: src/VX_elastic_buffer.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_elastic_buffer.sv:3:15
	parameter SIZE = 1;
	// Trace: src/VX_elastic_buffer.sv:4:15
	parameter OUT_REG = 0;
	// Trace: src/VX_elastic_buffer.sv:5:15
	parameter LUTRAM = 0;
	// Trace: src/VX_elastic_buffer.sv:7:5
	input wire clk;
	// Trace: src/VX_elastic_buffer.sv:8:5
	input wire reset;
	// Trace: src/VX_elastic_buffer.sv:9:5
	input wire valid_in;
	// Trace: src/VX_elastic_buffer.sv:10:5
	output wire ready_in;
	// Trace: src/VX_elastic_buffer.sv:11:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_elastic_buffer.sv:12:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_elastic_buffer.sv:13:5
	input wire ready_out;
	// Trace: src/VX_elastic_buffer.sv:14:5
	output wire valid_out;
	// Trace: src/VX_elastic_buffer.sv:16:5
	generate
		if (SIZE == 0) begin : g_passthru
			// Trace: src/VX_elastic_buffer.sv:17:9
			assign valid_out = valid_in;
			// Trace: src/VX_elastic_buffer.sv:18:9
			assign data_out = data_in;
			// Trace: src/VX_elastic_buffer.sv:19:9
			assign ready_in = ready_out;
		end
		else if (SIZE == 1) begin : g_eb1
			// Trace: src/VX_elastic_buffer.sv:21:9
			VX_pipe_buffer #(
				.DATAW(DATAW),
				.DEPTH((OUT_REG > 1 ? OUT_REG : 1))
			) pipe_buffer(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_in),
				.data_in(data_in),
				.ready_in(ready_in),
				.valid_out(valid_out),
				.data_out(data_out),
				.ready_out(ready_out)
			);
		end
		else if ((SIZE == 2) && (LUTRAM == 0)) begin : g_eb2
			// Trace: src/VX_elastic_buffer.sv:35:9
			wire valid_out_t;
			// Trace: src/VX_elastic_buffer.sv:36:9
			wire [DATAW - 1:0] data_out_t;
			// Trace: src/VX_elastic_buffer.sv:37:9
			wire ready_out_t;
			// Trace: src/VX_elastic_buffer.sv:38:9
			VX_stream_buffer #(
				.DATAW(DATAW),
				.OUT_REG(OUT_REG == 1)
			) stream_buffer(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_in),
				.data_in(data_in),
				.ready_in(ready_in),
				.valid_out(valid_out_t),
				.data_out(data_out_t),
				.ready_out(ready_out_t)
			);
			// Trace: src/VX_elastic_buffer.sv:51:9
			VX_pipe_buffer #(
				.DATAW(DATAW),
				.DEPTH((OUT_REG > 1 ? OUT_REG - 1 : 0))
			) out_buf(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_out_t),
				.data_in(data_out_t),
				.ready_in(ready_out_t),
				.valid_out(valid_out),
				.data_out(data_out),
				.ready_out(ready_out)
			);
		end
		else begin : g_ebN
			// Trace: src/VX_elastic_buffer.sv:65:9
			wire empty;
			wire full;
			// Trace: src/VX_elastic_buffer.sv:66:9
			wire [DATAW - 1:0] data_out_t;
			// Trace: src/VX_elastic_buffer.sv:67:9
			wire ready_out_t;
			// Trace: src/VX_elastic_buffer.sv:68:9
			wire valid_out_t = ~empty;
			// Trace: src/VX_elastic_buffer.sv:69:9
			wire push = valid_in && ready_in;
			// Trace: src/VX_elastic_buffer.sv:70:9
			wire pop = valid_out_t && ready_out_t;
			// Trace: src/VX_elastic_buffer.sv:71:9
			VX_fifo_queue #(
				.DATAW(DATAW),
				.DEPTH(SIZE),
				.OUT_REG(OUT_REG == 1),
				.LUTRAM(LUTRAM)
			) fifo_queue(
				.clk(clk),
				.reset(reset),
				.push(push),
				.pop(pop),
				.data_in(data_in),
				.data_out(data_out_t),
				.empty(empty),
				.full(full),
				.alm_empty(),
				.alm_full(),
				.size()
			);
			// Trace: src/VX_elastic_buffer.sv:89:9
			assign ready_in = ~full;
			// Trace: src/VX_elastic_buffer.sv:90:9
			VX_pipe_buffer #(
				.DATAW(DATAW),
				.DEPTH((OUT_REG > 1 ? OUT_REG - 1 : 0))
			) out_buf(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_out_t),
				.data_in(data_out_t),
				.ready_in(ready_out_t),
				.valid_out(valid_out),
				.data_out(data_out),
				.ready_out(ready_out)
			);
		end
	endgenerate
endmodule
module VX_allocator (
	clk,
	reset,
	acquire_en,
	acquire_addr,
	release_en,
	release_addr,
	empty,
	full
);
	// Trace: src/VX_allocator.sv:2:15
	parameter SIZE = 1;
	// Trace: src/VX_allocator.sv:3:15
	parameter ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
	// Trace: src/VX_allocator.sv:5:5
	input wire clk;
	// Trace: src/VX_allocator.sv:6:5
	input wire reset;
	// Trace: src/VX_allocator.sv:7:5
	input wire acquire_en;
	// Trace: src/VX_allocator.sv:8:5
	output wire [ADDRW - 1:0] acquire_addr;
	// Trace: src/VX_allocator.sv:9:5
	input wire release_en;
	// Trace: src/VX_allocator.sv:10:5
	input wire [ADDRW - 1:0] release_addr;
	// Trace: src/VX_allocator.sv:11:5
	output wire empty;
	// Trace: src/VX_allocator.sv:12:5
	output wire full;
	// Trace: src/VX_allocator.sv:14:5
	reg [SIZE - 1:0] free_slots;
	reg [SIZE - 1:0] free_slots_n;
	// Trace: src/VX_allocator.sv:15:5
	reg [ADDRW - 1:0] acquire_addr_r;
	// Trace: src/VX_allocator.sv:16:5
	reg empty_r;
	reg full_r;
	// Trace: src/VX_allocator.sv:17:5
	wire [ADDRW - 1:0] free_index;
	// Trace: src/VX_allocator.sv:18:5
	wire free_valid;
	// Trace: src/VX_allocator.sv:19:5
	always @(*) begin
		// Trace: src/VX_allocator.sv:20:9
		free_slots_n = free_slots;
		// Trace: src/VX_allocator.sv:21:9
		if (release_en)
			// Trace: src/VX_allocator.sv:22:13
			free_slots_n[release_addr] = 1;
		if (acquire_en)
			// Trace: src/VX_allocator.sv:25:13
			free_slots_n[acquire_addr_r] = 0;
	end
	// Trace: src/VX_allocator.sv:28:5
	VX_lzc #(
		.N(SIZE),
		.REVERSE(1)
	) free_slots_sel(
		.data_in(free_slots_n),
		.data_out(free_index),
		.valid_out(free_valid)
	);
	// Trace: src/VX_allocator.sv:36:5
	function automatic [ADDRW - 1:0] sv2v_cast_8BB5D;
		input reg [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D = inp;
	endfunction
	always @(posedge clk)
		// Trace: src/VX_allocator.sv:37:9
		if (reset) begin
			// Trace: src/VX_allocator.sv:38:13
			acquire_addr_r <= sv2v_cast_8BB5D(1'b0);
			// Trace: src/VX_allocator.sv:39:13
			free_slots <= {SIZE {1'b1}};
			// Trace: src/VX_allocator.sv:40:13
			empty_r <= 1'b1;
			// Trace: src/VX_allocator.sv:41:13
			full_r <= 1'b0;
		end
		else begin
			// Trace: src/VX_allocator.sv:43:13
			if (release_en)
				;
			if (acquire_en)
				;
			if (acquire_en || (release_en && full_r))
				// Trace: src/VX_allocator.sv:50:17
				acquire_addr_r <= free_index;
			// Trace: src/VX_allocator.sv:52:13
			free_slots <= free_slots_n;
			// Trace: src/VX_allocator.sv:53:13
			empty_r <= &free_slots_n;
			// Trace: src/VX_allocator.sv:54:13
			full_r <= ~free_valid;
		end
	// Trace: src/VX_allocator.sv:57:5
	assign acquire_addr = acquire_addr_r;
	// Trace: src/VX_allocator.sv:58:5
	assign empty = empty_r;
	// Trace: src/VX_allocator.sv:59:5
	assign full = full_r;
endmodule
// removed module with interface ports: VX_sfu_unit
// removed interface: VX_mem_bus_if
module VX_stream_arb (
	clk,
	reset,
	valid_in,
	data_in,
	ready_in,
	valid_out,
	data_out,
	ready_out,
	sel_out
);
	// Trace: src/VX_stream_arb.sv:2:15
	parameter NUM_INPUTS = 1;
	// Trace: src/VX_stream_arb.sv:3:15
	parameter NUM_OUTPUTS = 1;
	// Trace: src/VX_stream_arb.sv:4:15
	parameter DATAW = 1;
	// Trace: src/VX_stream_arb.sv:5:15
	parameter ARBITER = "R";
	// Trace: src/VX_stream_arb.sv:6:15
	parameter MAX_FANOUT = 8;
	// Trace: src/VX_stream_arb.sv:7:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_arb.sv:8:15
	parameter NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
	// Trace: src/VX_stream_arb.sv:9:15
	parameter SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
	// Trace: src/VX_stream_arb.sv:10:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: src/VX_stream_arb.sv:11:15
	parameter NUM_REQS_W = (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1);
	// Trace: src/VX_stream_arb.sv:13:5
	input wire clk;
	// Trace: src/VX_stream_arb.sv:14:5
	input wire reset;
	// Trace: src/VX_stream_arb.sv:15:5
	input wire [NUM_INPUTS - 1:0] valid_in;
	// Trace: src/VX_stream_arb.sv:16:5
	input wire [(NUM_INPUTS * DATAW) - 1:0] data_in;
	// Trace: src/VX_stream_arb.sv:17:5
	output wire [NUM_INPUTS - 1:0] ready_in;
	// Trace: src/VX_stream_arb.sv:18:5
	output wire [NUM_OUTPUTS - 1:0] valid_out;
	// Trace: src/VX_stream_arb.sv:19:5
	output wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out;
	// Trace: src/VX_stream_arb.sv:20:5
	input wire [NUM_OUTPUTS - 1:0] ready_out;
	// Trace: src/VX_stream_arb.sv:21:5
	output wire [(SEL_COUNT * NUM_REQS_W) - 1:0] sel_out;
	// Trace: src/VX_stream_arb.sv:23:5
	function automatic signed [NUM_REQS_W - 1:0] sv2v_cast_A9560_signed;
		input reg signed [NUM_REQS_W - 1:0] inp;
		sv2v_cast_A9560_signed = inp;
	endfunction
	generate
		if (NUM_INPUTS > NUM_OUTPUTS) begin : g_input_select
			if ((MAX_FANOUT != 0) && (NUM_REQS > (MAX_FANOUT + (MAX_FANOUT / 2)))) begin : g_fanout
				// Trace: src/VX_stream_arb.sv:25:13
				localparam NUM_SLICES = ((NUM_REQS + MAX_FANOUT) - 1) / MAX_FANOUT;
				// Trace: src/VX_stream_arb.sv:26:13
				localparam LOG_NUM_REQS2 = $clog2(MAX_FANOUT);
				// Trace: src/VX_stream_arb.sv:27:13
				localparam LOG_NUM_REQS3 = $clog2(NUM_SLICES);
				// Trace: src/VX_stream_arb.sv:28:13
				localparam DATAW2 = DATAW + LOG_NUM_REQS2;
				// Trace: src/VX_stream_arb.sv:29:13
				wire [(NUM_SLICES * NUM_OUTPUTS) - 1:0] valid_tmp;
				// Trace: src/VX_stream_arb.sv:30:13
				wire [((NUM_SLICES * NUM_OUTPUTS) * DATAW2) - 1:0] data_tmp;
				// Trace: src/VX_stream_arb.sv:31:13
				wire [(NUM_SLICES * NUM_OUTPUTS) - 1:0] ready_tmp;
				genvar _gv_s_2;
				for (_gv_s_2 = 0; _gv_s_2 < NUM_SLICES; _gv_s_2 = _gv_s_2 + 1) begin : g_slice_arbs
					localparam s = _gv_s_2;
					// Trace: src/VX_stream_arb.sv:33:17
					localparam SLICE_STRIDE = MAX_FANOUT * NUM_OUTPUTS;
					// Trace: src/VX_stream_arb.sv:34:17
					localparam SLICE_BEGIN = s * SLICE_STRIDE;
					// Trace: src/VX_stream_arb.sv:35:17
					localparam SLICE_END = ((SLICE_BEGIN + SLICE_STRIDE) < NUM_INPUTS ? SLICE_BEGIN + SLICE_STRIDE : NUM_INPUTS);
					// Trace: src/VX_stream_arb.sv:36:17
					localparam SLICE_SIZE = SLICE_END - SLICE_BEGIN;
					// Trace: src/VX_stream_arb.sv:37:17
					wire [(NUM_OUTPUTS * DATAW) - 1:0] data_tmp_u;
					// Trace: src/VX_stream_arb.sv:38:17
					wire [(NUM_OUTPUTS * LOG_NUM_REQS2) - 1:0] sel_tmp_u;
					// Trace: src/VX_stream_arb.sv:39:17
					VX_stream_arb #(
						.NUM_INPUTS(SLICE_SIZE),
						.NUM_OUTPUTS(NUM_OUTPUTS),
						.DATAW(DATAW),
						.ARBITER(ARBITER),
						.MAX_FANOUT(MAX_FANOUT),
						.OUT_BUF(3)
					) fanout_slice_arb(
						.clk(clk),
						.reset(reset),
						.valid_in(valid_in[SLICE_END - 1:SLICE_BEGIN]),
						.data_in(data_in[DATAW * (((SLICE_END - 1) >= SLICE_BEGIN ? SLICE_END - 1 : ((SLICE_END - 1) + ((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1)) - 1) - (((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1) - 1))+:DATAW * ((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1)]),
						.ready_in(ready_in[SLICE_END - 1:SLICE_BEGIN]),
						.valid_out(valid_tmp[s * NUM_OUTPUTS+:NUM_OUTPUTS]),
						.data_out(data_tmp_u),
						.ready_out(ready_tmp[s * NUM_OUTPUTS+:NUM_OUTPUTS]),
						.sel_out(sel_tmp_u)
					);
					genvar _gv_o_1;
					for (_gv_o_1 = 0; _gv_o_1 < NUM_OUTPUTS; _gv_o_1 = _gv_o_1 + 1) begin : g_data_tmp
						localparam o = _gv_o_1;
						// Trace: src/VX_stream_arb.sv:58:21
						assign data_tmp[((s * NUM_OUTPUTS) + o) * DATAW2+:DATAW2] = {data_tmp_u[o * DATAW+:DATAW], sel_tmp_u[o * LOG_NUM_REQS2+:LOG_NUM_REQS2]};
					end
				end
				// Trace: src/VX_stream_arb.sv:61:13
				wire [(NUM_OUTPUTS * DATAW2) - 1:0] data_out_u;
				// Trace: src/VX_stream_arb.sv:62:13
				wire [(NUM_OUTPUTS * LOG_NUM_REQS3) - 1:0] sel_out_u;
				// Trace: src/VX_stream_arb.sv:63:13
				VX_stream_arb #(
					.NUM_INPUTS(NUM_SLICES * NUM_OUTPUTS),
					.NUM_OUTPUTS(NUM_OUTPUTS),
					.DATAW(DATAW2),
					.ARBITER(ARBITER),
					.MAX_FANOUT(MAX_FANOUT),
					.OUT_BUF(OUT_BUF)
				) fanout_join_arb(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_tmp),
					.ready_in(ready_tmp),
					.data_in(data_tmp),
					.data_out(data_out_u),
					.sel_out(sel_out_u),
					.valid_out(valid_out),
					.ready_out(ready_out)
				);
				genvar _gv_o_2;
				for (_gv_o_2 = 0; _gv_o_2 < NUM_OUTPUTS; _gv_o_2 = _gv_o_2 + 1) begin : g_data_out
					localparam o = _gv_o_2;
					// Trace: src/VX_stream_arb.sv:82:17
					assign sel_out[o * NUM_REQS_W+:NUM_REQS_W] = {sel_out_u[o * LOG_NUM_REQS3+:LOG_NUM_REQS3], data_out_u[(o * DATAW2) + (LOG_NUM_REQS2 - 1)-:LOG_NUM_REQS2]};
					// Trace: src/VX_stream_arb.sv:83:17
					assign data_out[o * DATAW+:DATAW] = data_out_u[(o * DATAW2) + ((DATAW2 - 1) >= LOG_NUM_REQS2 ? DATAW2 - 1 : ((DATAW2 - 1) + ((DATAW2 - 1) >= LOG_NUM_REQS2 ? ((DATAW2 - 1) - LOG_NUM_REQS2) + 1 : (LOG_NUM_REQS2 - (DATAW2 - 1)) + 1)) - 1)-:((DATAW2 - 1) >= LOG_NUM_REQS2 ? ((DATAW2 - 1) - LOG_NUM_REQS2) + 1 : (LOG_NUM_REQS2 - (DATAW2 - 1)) + 1)];
				end
			end
			else begin : g_arbiter
				// Trace: src/VX_stream_arb.sv:86:13
				wire [NUM_REQS - 1:0] arb_requests;
				// Trace: src/VX_stream_arb.sv:87:13
				wire arb_valid;
				// Trace: src/VX_stream_arb.sv:88:13
				wire [NUM_REQS_W - 1:0] arb_index;
				// Trace: src/VX_stream_arb.sv:89:13
				wire [NUM_REQS - 1:0] arb_onehot;
				// Trace: src/VX_stream_arb.sv:90:13
				wire arb_ready;
				genvar _gv_r_7;
				for (_gv_r_7 = 0; _gv_r_7 < NUM_REQS; _gv_r_7 = _gv_r_7 + 1) begin : g_requests
					localparam r = _gv_r_7;
					// Trace: src/VX_stream_arb.sv:92:17
					wire [NUM_OUTPUTS - 1:0] requests;
					genvar _gv_o_3;
					for (_gv_o_3 = 0; _gv_o_3 < NUM_OUTPUTS; _gv_o_3 = _gv_o_3 + 1) begin : g_o
						localparam o = _gv_o_3;
						// Trace: src/VX_stream_arb.sv:94:21
						localparam i = (r * NUM_OUTPUTS) + o;
						// Trace: src/VX_stream_arb.sv:95:21
						assign requests[o] = valid_in[i];
					end
					// Trace: src/VX_stream_arb.sv:97:17
					assign arb_requests[r] = |requests;
				end
				// Trace: src/VX_stream_arb.sv:99:13
				VX_generic_arbiter #(
					.NUM_REQS(NUM_REQS),
					.TYPE(ARBITER)
				) arbiter(
					.clk(clk),
					.reset(reset),
					.requests(arb_requests),
					.grant_valid(arb_valid),
					.grant_index(arb_index),
					.grant_onehot(arb_onehot),
					.grant_ready(arb_ready)
				);
				// Trace: src/VX_stream_arb.sv:111:13
				wire [NUM_OUTPUTS - 1:0] valid_out_w;
				// Trace: src/VX_stream_arb.sv:112:13
				wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out_w;
				// Trace: src/VX_stream_arb.sv:113:13
				wire [NUM_OUTPUTS - 1:0] ready_out_w;
				genvar _gv_o_4;
				for (_gv_o_4 = 0; _gv_o_4 < NUM_OUTPUTS; _gv_o_4 = _gv_o_4 + 1) begin : g_data_out_w
					localparam o = _gv_o_4;
					// Trace: src/VX_stream_arb.sv:115:17
					wire [NUM_REQS - 1:0] valid_in_w;
					// Trace: src/VX_stream_arb.sv:116:17
					wire [(NUM_REQS * DATAW) - 1:0] data_in_w;
					genvar _gv_r_8;
					for (_gv_r_8 = 0; _gv_r_8 < NUM_REQS; _gv_r_8 = _gv_r_8 + 1) begin : g_r
						localparam r = _gv_r_8;
						// Trace: src/VX_stream_arb.sv:118:21
						localparam i = (r * NUM_OUTPUTS) + o;
						if (r < NUM_INPUTS) begin : g_valid
							// Trace: src/VX_stream_arb.sv:120:25
							assign valid_in_w[r] = valid_in[i];
							// Trace: src/VX_stream_arb.sv:121:25
							assign data_in_w[r * DATAW+:DATAW] = data_in[i * DATAW+:DATAW];
						end
						else begin : g_padding
							// Trace: src/VX_stream_arb.sv:123:25
							assign valid_in_w[r] = 0;
							// Trace: src/VX_stream_arb.sv:124:25
							assign data_in_w[r * DATAW+:DATAW] = 1'sb0;
						end
					end
					// Trace: src/VX_stream_arb.sv:127:17
					assign valid_out_w[o] = (NUM_OUTPUTS == 1 ? arb_valid : |(valid_in_w & arb_onehot));
					// Trace: src/VX_stream_arb.sv:128:17
					assign data_out_w[o * DATAW+:DATAW] = data_in_w[arb_index * DATAW+:DATAW];
				end
				genvar _gv_i_158;
				for (_gv_i_158 = 0; _gv_i_158 < NUM_INPUTS; _gv_i_158 = _gv_i_158 + 1) begin : g_ready_in
					localparam i = _gv_i_158;
					// Trace: src/VX_stream_arb.sv:131:17
					localparam o = i % NUM_OUTPUTS;
					// Trace: src/VX_stream_arb.sv:132:17
					localparam r = i / NUM_OUTPUTS;
					// Trace: src/VX_stream_arb.sv:133:17
					assign ready_in[i] = ready_out_w[o] && arb_onehot[r];
				end
				// Trace: src/VX_stream_arb.sv:135:13
				assign arb_ready = |ready_out_w;
				genvar _gv_o_5;
				for (_gv_o_5 = 0; _gv_o_5 < NUM_OUTPUTS; _gv_o_5 = _gv_o_5 + 1) begin : g_out_buf
					localparam o = _gv_o_5;
					// Trace: src/VX_stream_arb.sv:137:17
					VX_elastic_buffer #(
						.DATAW(LOG_NUM_REQS + DATAW),
						.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
						.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
						.LUTRAM((OUT_BUF & 8) != 0)
					) out_buf(
						.clk(clk),
						.reset(reset),
						.valid_in(valid_out_w[o]),
						.ready_in(ready_out_w[o]),
						.data_in({arb_index, data_out_w[o * DATAW+:DATAW]}),
						.data_out({sel_out[o * NUM_REQS_W+:NUM_REQS_W], data_out[o * DATAW+:DATAW]}),
						.valid_out(valid_out[o]),
						.ready_out(ready_out[o])
					);
				end
			end
		end
		else if (NUM_INPUTS < NUM_OUTPUTS) begin : g_output_select
			if ((MAX_FANOUT != 0) && (NUM_REQS > (MAX_FANOUT + (MAX_FANOUT / 2)))) begin : g_fanout
				// Trace: src/VX_stream_arb.sv:156:13
				localparam NUM_SLICES = ((NUM_REQS + MAX_FANOUT) - 1) / MAX_FANOUT;
				// Trace: src/VX_stream_arb.sv:157:13
				localparam LOG_NUM_REQS2 = $clog2(MAX_FANOUT);
				// Trace: src/VX_stream_arb.sv:158:13
				localparam LOG_NUM_REQS3 = $clog2(NUM_SLICES);
				// Trace: src/VX_stream_arb.sv:159:13
				wire [(NUM_SLICES * NUM_INPUTS) - 1:0] valid_tmp;
				// Trace: src/VX_stream_arb.sv:160:13
				wire [((NUM_SLICES * NUM_INPUTS) * DATAW) - 1:0] data_tmp;
				// Trace: src/VX_stream_arb.sv:161:13
				wire [(NUM_SLICES * NUM_INPUTS) - 1:0] ready_tmp;
				// Trace: src/VX_stream_arb.sv:162:13
				wire [(NUM_INPUTS * LOG_NUM_REQS3) - 1:0] sel_tmp;
				// Trace: src/VX_stream_arb.sv:163:13
				VX_stream_arb #(
					.NUM_INPUTS(NUM_INPUTS),
					.NUM_OUTPUTS(NUM_SLICES * NUM_INPUTS),
					.DATAW(DATAW),
					.ARBITER(ARBITER),
					.MAX_FANOUT(MAX_FANOUT),
					.OUT_BUF(3)
				) fanout_fork_arb(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_in),
					.ready_in(ready_in),
					.data_in(data_in),
					.data_out(data_tmp),
					.valid_out(valid_tmp),
					.ready_out(ready_tmp),
					.sel_out(sel_tmp)
				);
				// Trace: src/VX_stream_arb.sv:181:13
				wire [((NUM_SLICES * NUM_INPUTS) * LOG_NUM_REQS2) - 1:0] sel_out_w;
				genvar _gv_s_3;
				for (_gv_s_3 = 0; _gv_s_3 < NUM_SLICES; _gv_s_3 = _gv_s_3 + 1) begin : g_slice_arbs
					localparam s = _gv_s_3;
					// Trace: src/VX_stream_arb.sv:183:17
					localparam SLICE_STRIDE = MAX_FANOUT * NUM_INPUTS;
					// Trace: src/VX_stream_arb.sv:184:17
					localparam SLICE_BEGIN = s * SLICE_STRIDE;
					// Trace: src/VX_stream_arb.sv:185:17
					localparam SLICE_END = ((SLICE_BEGIN + SLICE_STRIDE) < NUM_OUTPUTS ? SLICE_BEGIN + SLICE_STRIDE : NUM_OUTPUTS);
					// Trace: src/VX_stream_arb.sv:186:17
					localparam SLICE_SIZE = SLICE_END - SLICE_BEGIN;
					// Trace: src/VX_stream_arb.sv:187:17
					wire [(NUM_INPUTS * LOG_NUM_REQS2) - 1:0] sel_out_u;
					// Trace: src/VX_stream_arb.sv:188:17
					VX_stream_arb #(
						.NUM_INPUTS(NUM_INPUTS),
						.NUM_OUTPUTS(SLICE_SIZE),
						.DATAW(DATAW),
						.ARBITER(ARBITER),
						.MAX_FANOUT(MAX_FANOUT),
						.OUT_BUF(OUT_BUF)
					) fanout_slice_arb(
						.clk(clk),
						.reset(reset),
						.valid_in(valid_tmp[s * NUM_INPUTS+:NUM_INPUTS]),
						.ready_in(ready_tmp[s * NUM_INPUTS+:NUM_INPUTS]),
						.data_in(data_tmp[DATAW * (s * NUM_INPUTS)+:DATAW * NUM_INPUTS]),
						.data_out(data_out[DATAW * (((SLICE_END - 1) >= SLICE_BEGIN ? SLICE_END - 1 : ((SLICE_END - 1) + ((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1)) - 1) - (((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1) - 1))+:DATAW * ((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1)]),
						.valid_out(valid_out[SLICE_END - 1:SLICE_BEGIN]),
						.ready_out(ready_out[SLICE_END - 1:SLICE_BEGIN]),
						.sel_out(sel_out_w[LOG_NUM_REQS2 * (s * NUM_INPUTS)+:LOG_NUM_REQS2 * NUM_INPUTS])
					);
				end
				genvar _gv_i_159;
				for (_gv_i_159 = 0; _gv_i_159 < NUM_INPUTS; _gv_i_159 = _gv_i_159 + 1) begin : g_sel_out
					localparam i = _gv_i_159;
					// Trace: src/VX_stream_arb.sv:208:17
					assign sel_out[i * NUM_REQS_W+:NUM_REQS_W] = {sel_tmp[i * LOG_NUM_REQS3+:LOG_NUM_REQS3], sel_out_w[((sel_tmp[i * LOG_NUM_REQS3+:LOG_NUM_REQS3] * NUM_INPUTS) + i) * LOG_NUM_REQS2+:LOG_NUM_REQS2]};
				end
			end
			else begin : g_arbiter
				// Trace: src/VX_stream_arb.sv:211:13
				wire [NUM_REQS - 1:0] arb_requests;
				// Trace: src/VX_stream_arb.sv:212:13
				wire arb_valid;
				// Trace: src/VX_stream_arb.sv:213:13
				wire [NUM_REQS_W - 1:0] arb_index;
				// Trace: src/VX_stream_arb.sv:214:13
				wire [NUM_REQS - 1:0] arb_onehot;
				// Trace: src/VX_stream_arb.sv:215:13
				wire arb_ready;
				genvar _gv_r_9;
				for (_gv_r_9 = 0; _gv_r_9 < NUM_REQS; _gv_r_9 = _gv_r_9 + 1) begin : g_requests
					localparam r = _gv_r_9;
					// Trace: src/VX_stream_arb.sv:217:17
					wire [NUM_INPUTS - 1:0] requests;
					genvar _gv_i_160;
					for (_gv_i_160 = 0; _gv_i_160 < NUM_INPUTS; _gv_i_160 = _gv_i_160 + 1) begin : g_i
						localparam i = _gv_i_160;
						// Trace: src/VX_stream_arb.sv:219:21
						localparam o = (r * NUM_INPUTS) + i;
						// Trace: src/VX_stream_arb.sv:220:21
						assign requests[i] = ready_out[o];
					end
					// Trace: src/VX_stream_arb.sv:222:17
					assign arb_requests[r] = |requests;
				end
				// Trace: src/VX_stream_arb.sv:224:13
				VX_generic_arbiter #(
					.NUM_REQS(NUM_REQS),
					.TYPE(ARBITER)
				) arbiter(
					.clk(clk),
					.reset(reset),
					.requests(arb_requests),
					.grant_valid(arb_valid),
					.grant_index(arb_index),
					.grant_onehot(arb_onehot),
					.grant_ready(arb_ready)
				);
				// Trace: src/VX_stream_arb.sv:236:13
				wire [NUM_OUTPUTS - 1:0] valid_out_w;
				// Trace: src/VX_stream_arb.sv:237:13
				wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out_w;
				// Trace: src/VX_stream_arb.sv:238:13
				wire [NUM_OUTPUTS - 1:0] ready_out_w;
				genvar _gv_o_6;
				for (_gv_o_6 = 0; _gv_o_6 < NUM_OUTPUTS; _gv_o_6 = _gv_o_6 + 1) begin : g_data_out_w
					localparam o = _gv_o_6;
					// Trace: src/VX_stream_arb.sv:240:17
					localparam i = o % NUM_INPUTS;
					// Trace: src/VX_stream_arb.sv:241:17
					localparam r = o / NUM_INPUTS;
					// Trace: src/VX_stream_arb.sv:242:17
					assign valid_out_w[o] = valid_in[i] && arb_onehot[r];
					// Trace: src/VX_stream_arb.sv:243:17
					assign data_out_w[o * DATAW+:DATAW] = data_in[i * DATAW+:DATAW];
				end
				genvar _gv_i_161;
				for (_gv_i_161 = 0; _gv_i_161 < NUM_INPUTS; _gv_i_161 = _gv_i_161 + 1) begin : g_ready_in
					localparam i = _gv_i_161;
					// Trace: src/VX_stream_arb.sv:246:17
					wire [NUM_REQS - 1:0] ready_out_s;
					genvar _gv_r_10;
					for (_gv_r_10 = 0; _gv_r_10 < NUM_REQS; _gv_r_10 = _gv_r_10 + 1) begin : g_r
						localparam r = _gv_r_10;
						// Trace: src/VX_stream_arb.sv:248:21
						localparam o = (r * NUM_INPUTS) + i;
						// Trace: src/VX_stream_arb.sv:249:21
						assign ready_out_s[r] = ready_out_w[o];
					end
					// Trace: src/VX_stream_arb.sv:251:17
					assign ready_in[i] = (NUM_INPUTS == 1 ? arb_valid : |(ready_out_s & arb_onehot));
				end
				// Trace: src/VX_stream_arb.sv:253:13
				assign arb_ready = |valid_in;
				genvar _gv_o_7;
				for (_gv_o_7 = 0; _gv_o_7 < NUM_OUTPUTS; _gv_o_7 = _gv_o_7 + 1) begin : g_out_buf
					localparam o = _gv_o_7;
					// Trace: src/VX_stream_arb.sv:255:17
					VX_elastic_buffer #(
						.DATAW(DATAW),
						.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
						.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
						.LUTRAM((OUT_BUF & 8) != 0)
					) out_buf(
						.clk(clk),
						.reset(reset),
						.valid_in(valid_out_w[o]),
						.ready_in(ready_out_w[o]),
						.data_in(data_out_w[o * DATAW+:DATAW]),
						.data_out(data_out[o * DATAW+:DATAW]),
						.valid_out(valid_out[o]),
						.ready_out(ready_out[o])
					);
				end
				genvar _gv_i_162;
				for (_gv_i_162 = 0; _gv_i_162 < NUM_INPUTS; _gv_i_162 = _gv_i_162 + 1) begin : g_sel_out
					localparam i = _gv_i_162;
					// Trace: src/VX_stream_arb.sv:272:17
					assign sel_out[i * NUM_REQS_W+:NUM_REQS_W] = arb_index;
				end
			end
		end
		else begin : g_passthru
			genvar _gv_o_8;
			for (_gv_o_8 = 0; _gv_o_8 < NUM_OUTPUTS; _gv_o_8 = _gv_o_8 + 1) begin : g_out_buf
				localparam o = _gv_o_8;
				// Trace: src/VX_stream_arb.sv:277:13
				VX_elastic_buffer #(
					.DATAW(DATAW),
					.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
					.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
					.LUTRAM((OUT_BUF & 8) != 0)
				) out_buf(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_in[o]),
					.ready_in(ready_in[o]),
					.data_in(data_in[o * DATAW+:DATAW]),
					.data_out(data_out[o * DATAW+:DATAW]),
					.valid_out(valid_out[o]),
					.ready_out(ready_out[o])
				);
				// Trace: src/VX_stream_arb.sv:292:13
				assign sel_out[o * NUM_REQS_W+:NUM_REQS_W] = sv2v_cast_A9560_signed(0);
			end
		end
	endgenerate
endmodule
module VX_bits_remove (
	data_in,
	sel_out,
	data_out
);
	// Trace: src/VX_bits_remove.sv:2:15
	parameter N = 2;
	// Trace: src/VX_bits_remove.sv:3:15
	parameter S = 1;
	// Trace: src/VX_bits_remove.sv:4:15
	parameter POS = 0;
	// Trace: src/VX_bits_remove.sv:6:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_bits_remove.sv:7:5
	output wire [(S > 0 ? S : 1) - 1:0] sel_out;
	// Trace: src/VX_bits_remove.sv:8:5
	output wire [(N - S) - 1:0] data_out;
	// Trace: src/VX_bits_remove.sv:10:5
	generate
		if (S == 0) begin : g_passthru
			// Trace: src/VX_bits_remove.sv:11:9
			assign sel_out = 0;
			// Trace: src/VX_bits_remove.sv:12:9
			assign data_out = data_in;
		end
		else if (POS == 0) begin : g_pos_0
			// Trace: src/VX_bits_remove.sv:14:9
			assign sel_out = data_in[0+:S];
			// Trace: src/VX_bits_remove.sv:15:9
			assign data_out = data_in[N - 1:S];
		end
		else if ((POS + S) == N) begin : g_pos_N
			// Trace: src/VX_bits_remove.sv:17:9
			assign sel_out = data_in[POS+:S];
			// Trace: src/VX_bits_remove.sv:18:9
			assign data_out = data_in[POS - 1:0];
		end
		else begin : g_pos
			// Trace: src/VX_bits_remove.sv:20:9
			assign sel_out = data_in[POS+:S];
			// Trace: src/VX_bits_remove.sv:21:9
			assign data_out = {data_in[N - 1:POS + S], data_in[POS - 1:0]};
		end
	endgenerate
endmodule
// removed module with interface ports: VX_execute
// removed module with interface ports: VX_gbar_arb
module VX_popcount63 (
	data_in,
	data_out
);
	// Trace: src/VX_popcount.sv:2:5
	input wire [5:0] data_in;
	// Trace: src/VX_popcount.sv:3:5
	output wire [2:0] data_out;
	// Trace: src/VX_popcount.sv:5:5
	reg [2:0] sum;
	// Trace: src/VX_popcount.sv:6:5
	always @(*)
		// Trace: src/VX_popcount.sv:7:9
		case (data_in)
			6'd0:
				// Trace: src/VX_popcount.sv:8:16
				sum = 3'd0;
			6'd1:
				// Trace: src/VX_popcount.sv:8:34
				sum = 3'd1;
			6'd2:
				// Trace: src/VX_popcount.sv:8:52
				sum = 3'd1;
			6'd3:
				// Trace: src/VX_popcount.sv:8:70
				sum = 3'd2;
			6'd4:
				// Trace: src/VX_popcount.sv:9:16
				sum = 3'd1;
			6'd5:
				// Trace: src/VX_popcount.sv:9:34
				sum = 3'd2;
			6'd6:
				// Trace: src/VX_popcount.sv:9:52
				sum = 3'd2;
			6'd7:
				// Trace: src/VX_popcount.sv:9:70
				sum = 3'd3;
			6'd8:
				// Trace: src/VX_popcount.sv:10:16
				sum = 3'd1;
			6'd9:
				// Trace: src/VX_popcount.sv:10:34
				sum = 3'd2;
			6'd10:
				// Trace: src/VX_popcount.sv:10:52
				sum = 3'd2;
			6'd11:
				// Trace: src/VX_popcount.sv:10:70
				sum = 3'd3;
			6'd12:
				// Trace: src/VX_popcount.sv:11:16
				sum = 3'd2;
			6'd13:
				// Trace: src/VX_popcount.sv:11:34
				sum = 3'd3;
			6'd14:
				// Trace: src/VX_popcount.sv:11:52
				sum = 3'd3;
			6'd15:
				// Trace: src/VX_popcount.sv:11:70
				sum = 3'd4;
			6'd16:
				// Trace: src/VX_popcount.sv:12:16
				sum = 3'd1;
			6'd17:
				// Trace: src/VX_popcount.sv:12:34
				sum = 3'd2;
			6'd18:
				// Trace: src/VX_popcount.sv:12:52
				sum = 3'd2;
			6'd19:
				// Trace: src/VX_popcount.sv:12:70
				sum = 3'd3;
			6'd20:
				// Trace: src/VX_popcount.sv:13:16
				sum = 3'd2;
			6'd21:
				// Trace: src/VX_popcount.sv:13:34
				sum = 3'd3;
			6'd22:
				// Trace: src/VX_popcount.sv:13:52
				sum = 3'd3;
			6'd23:
				// Trace: src/VX_popcount.sv:13:70
				sum = 3'd4;
			6'd24:
				// Trace: src/VX_popcount.sv:14:16
				sum = 3'd2;
			6'd25:
				// Trace: src/VX_popcount.sv:14:34
				sum = 3'd3;
			6'd26:
				// Trace: src/VX_popcount.sv:14:52
				sum = 3'd3;
			6'd27:
				// Trace: src/VX_popcount.sv:14:70
				sum = 3'd4;
			6'd28:
				// Trace: src/VX_popcount.sv:15:16
				sum = 3'd3;
			6'd29:
				// Trace: src/VX_popcount.sv:15:34
				sum = 3'd4;
			6'd30:
				// Trace: src/VX_popcount.sv:15:52
				sum = 3'd4;
			6'd31:
				// Trace: src/VX_popcount.sv:15:70
				sum = 3'd5;
			6'd32:
				// Trace: src/VX_popcount.sv:16:16
				sum = 3'd1;
			6'd33:
				// Trace: src/VX_popcount.sv:16:34
				sum = 3'd2;
			6'd34:
				// Trace: src/VX_popcount.sv:16:52
				sum = 3'd2;
			6'd35:
				// Trace: src/VX_popcount.sv:16:70
				sum = 3'd3;
			6'd36:
				// Trace: src/VX_popcount.sv:17:16
				sum = 3'd2;
			6'd37:
				// Trace: src/VX_popcount.sv:17:34
				sum = 3'd3;
			6'd38:
				// Trace: src/VX_popcount.sv:17:52
				sum = 3'd3;
			6'd39:
				// Trace: src/VX_popcount.sv:17:70
				sum = 3'd4;
			6'd40:
				// Trace: src/VX_popcount.sv:18:16
				sum = 3'd2;
			6'd41:
				// Trace: src/VX_popcount.sv:18:34
				sum = 3'd3;
			6'd42:
				// Trace: src/VX_popcount.sv:18:52
				sum = 3'd3;
			6'd43:
				// Trace: src/VX_popcount.sv:18:70
				sum = 3'd4;
			6'd44:
				// Trace: src/VX_popcount.sv:19:16
				sum = 3'd3;
			6'd45:
				// Trace: src/VX_popcount.sv:19:34
				sum = 3'd4;
			6'd46:
				// Trace: src/VX_popcount.sv:19:52
				sum = 3'd4;
			6'd47:
				// Trace: src/VX_popcount.sv:19:70
				sum = 3'd5;
			6'd48:
				// Trace: src/VX_popcount.sv:20:16
				sum = 3'd2;
			6'd49:
				// Trace: src/VX_popcount.sv:20:34
				sum = 3'd3;
			6'd50:
				// Trace: src/VX_popcount.sv:20:52
				sum = 3'd3;
			6'd51:
				// Trace: src/VX_popcount.sv:20:70
				sum = 3'd4;
			6'd52:
				// Trace: src/VX_popcount.sv:21:16
				sum = 3'd3;
			6'd53:
				// Trace: src/VX_popcount.sv:21:34
				sum = 3'd4;
			6'd54:
				// Trace: src/VX_popcount.sv:21:52
				sum = 3'd4;
			6'd55:
				// Trace: src/VX_popcount.sv:21:70
				sum = 3'd5;
			6'd56:
				// Trace: src/VX_popcount.sv:22:16
				sum = 3'd3;
			6'd57:
				// Trace: src/VX_popcount.sv:22:34
				sum = 3'd4;
			6'd58:
				// Trace: src/VX_popcount.sv:22:52
				sum = 3'd4;
			6'd59:
				// Trace: src/VX_popcount.sv:22:70
				sum = 3'd5;
			6'd60:
				// Trace: src/VX_popcount.sv:23:16
				sum = 3'd4;
			6'd61:
				// Trace: src/VX_popcount.sv:23:34
				sum = 3'd5;
			6'd62:
				// Trace: src/VX_popcount.sv:23:52
				sum = 3'd5;
			6'd63:
				// Trace: src/VX_popcount.sv:23:70
				sum = 3'd6;
		endcase
	// Trace: src/VX_popcount.sv:26:5
	assign data_out = sum;
endmodule
module VX_popcount32 (
	data_in,
	data_out
);
	// Trace: src/VX_popcount.sv:29:5
	input wire [2:0] data_in;
	// Trace: src/VX_popcount.sv:30:5
	output wire [1:0] data_out;
	// Trace: src/VX_popcount.sv:32:5
	reg [1:0] sum;
	// Trace: src/VX_popcount.sv:33:5
	always @(*)
		// Trace: src/VX_popcount.sv:34:9
		case (data_in)
			3'd0:
				// Trace: src/VX_popcount.sv:35:15
				sum = 2'd0;
			3'd1:
				// Trace: src/VX_popcount.sv:35:33
				sum = 2'd1;
			3'd2:
				// Trace: src/VX_popcount.sv:35:51
				sum = 2'd1;
			3'd3:
				// Trace: src/VX_popcount.sv:35:69
				sum = 2'd2;
			3'd4:
				// Trace: src/VX_popcount.sv:36:15
				sum = 2'd1;
			3'd5:
				// Trace: src/VX_popcount.sv:36:33
				sum = 2'd2;
			3'd6:
				// Trace: src/VX_popcount.sv:36:51
				sum = 2'd2;
			3'd7:
				// Trace: src/VX_popcount.sv:36:69
				sum = 2'd3;
		endcase
	// Trace: src/VX_popcount.sv:39:5
	assign data_out = sum;
endmodule
module VX_sum33 (
	data_in1,
	data_in2,
	data_out
);
	// Trace: src/VX_popcount.sv:42:5
	input wire [2:0] data_in1;
	// Trace: src/VX_popcount.sv:43:5
	input wire [2:0] data_in2;
	// Trace: src/VX_popcount.sv:44:5
	output wire [3:0] data_out;
	// Trace: src/VX_popcount.sv:46:5
	reg [3:0] sum;
	// Trace: src/VX_popcount.sv:47:5
	always @(*)
		// Trace: src/VX_popcount.sv:48:9
		case ({data_in1, data_in2})
			6'd0:
				// Trace: src/VX_popcount.sv:49:16
				sum = 4'd0;
			6'd1:
				// Trace: src/VX_popcount.sv:49:34
				sum = 4'd1;
			6'd2:
				// Trace: src/VX_popcount.sv:49:52
				sum = 4'd2;
			6'd3:
				// Trace: src/VX_popcount.sv:49:70
				sum = 4'd3;
			6'd4:
				// Trace: src/VX_popcount.sv:50:16
				sum = 4'd4;
			6'd5:
				// Trace: src/VX_popcount.sv:50:34
				sum = 4'd5;
			6'd6:
				// Trace: src/VX_popcount.sv:50:52
				sum = 4'd6;
			6'd7:
				// Trace: src/VX_popcount.sv:50:70
				sum = 4'd7;
			6'd8:
				// Trace: src/VX_popcount.sv:51:16
				sum = 4'd1;
			6'd9:
				// Trace: src/VX_popcount.sv:51:34
				sum = 4'd2;
			6'd10:
				// Trace: src/VX_popcount.sv:51:52
				sum = 4'd3;
			6'd11:
				// Trace: src/VX_popcount.sv:51:70
				sum = 4'd4;
			6'd12:
				// Trace: src/VX_popcount.sv:52:16
				sum = 4'd5;
			6'd13:
				// Trace: src/VX_popcount.sv:52:34
				sum = 4'd6;
			6'd14:
				// Trace: src/VX_popcount.sv:52:52
				sum = 4'd7;
			6'd15:
				// Trace: src/VX_popcount.sv:52:70
				sum = 4'd8;
			6'd16:
				// Trace: src/VX_popcount.sv:53:16
				sum = 4'd2;
			6'd17:
				// Trace: src/VX_popcount.sv:53:34
				sum = 4'd3;
			6'd18:
				// Trace: src/VX_popcount.sv:53:52
				sum = 4'd4;
			6'd19:
				// Trace: src/VX_popcount.sv:53:70
				sum = 4'd5;
			6'd20:
				// Trace: src/VX_popcount.sv:54:16
				sum = 4'd6;
			6'd21:
				// Trace: src/VX_popcount.sv:54:34
				sum = 4'd7;
			6'd22:
				// Trace: src/VX_popcount.sv:54:52
				sum = 4'd8;
			6'd23:
				// Trace: src/VX_popcount.sv:54:70
				sum = 4'd9;
			6'd24:
				// Trace: src/VX_popcount.sv:55:16
				sum = 4'd3;
			6'd25:
				// Trace: src/VX_popcount.sv:55:34
				sum = 4'd4;
			6'd26:
				// Trace: src/VX_popcount.sv:55:52
				sum = 4'd5;
			6'd27:
				// Trace: src/VX_popcount.sv:55:70
				sum = 4'd6;
			6'd28:
				// Trace: src/VX_popcount.sv:56:16
				sum = 4'd7;
			6'd29:
				// Trace: src/VX_popcount.sv:56:34
				sum = 4'd8;
			6'd30:
				// Trace: src/VX_popcount.sv:56:52
				sum = 4'd9;
			6'd31:
				// Trace: src/VX_popcount.sv:56:70
				sum = 4'd10;
			6'd32:
				// Trace: src/VX_popcount.sv:57:16
				sum = 4'd4;
			6'd33:
				// Trace: src/VX_popcount.sv:57:34
				sum = 4'd5;
			6'd34:
				// Trace: src/VX_popcount.sv:57:52
				sum = 4'd6;
			6'd35:
				// Trace: src/VX_popcount.sv:57:70
				sum = 4'd7;
			6'd36:
				// Trace: src/VX_popcount.sv:58:16
				sum = 4'd8;
			6'd37:
				// Trace: src/VX_popcount.sv:58:34
				sum = 4'd9;
			6'd38:
				// Trace: src/VX_popcount.sv:58:52
				sum = 4'd10;
			6'd39:
				// Trace: src/VX_popcount.sv:58:70
				sum = 4'd11;
			6'd40:
				// Trace: src/VX_popcount.sv:59:16
				sum = 4'd5;
			6'd41:
				// Trace: src/VX_popcount.sv:59:34
				sum = 4'd6;
			6'd42:
				// Trace: src/VX_popcount.sv:59:52
				sum = 4'd7;
			6'd43:
				// Trace: src/VX_popcount.sv:59:70
				sum = 4'd8;
			6'd44:
				// Trace: src/VX_popcount.sv:60:16
				sum = 4'd9;
			6'd45:
				// Trace: src/VX_popcount.sv:60:34
				sum = 4'd10;
			6'd46:
				// Trace: src/VX_popcount.sv:60:52
				sum = 4'd11;
			6'd47:
				// Trace: src/VX_popcount.sv:60:70
				sum = 4'd12;
			6'd48:
				// Trace: src/VX_popcount.sv:61:16
				sum = 4'd6;
			6'd49:
				// Trace: src/VX_popcount.sv:61:34
				sum = 4'd7;
			6'd50:
				// Trace: src/VX_popcount.sv:61:52
				sum = 4'd8;
			6'd51:
				// Trace: src/VX_popcount.sv:61:70
				sum = 4'd9;
			6'd52:
				// Trace: src/VX_popcount.sv:62:16
				sum = 4'd10;
			6'd53:
				// Trace: src/VX_popcount.sv:62:34
				sum = 4'd11;
			6'd54:
				// Trace: src/VX_popcount.sv:62:52
				sum = 4'd12;
			6'd55:
				// Trace: src/VX_popcount.sv:62:70
				sum = 4'd13;
			6'd56:
				// Trace: src/VX_popcount.sv:63:16
				sum = 4'd7;
			6'd57:
				// Trace: src/VX_popcount.sv:63:34
				sum = 4'd8;
			6'd58:
				// Trace: src/VX_popcount.sv:63:52
				sum = 4'd9;
			6'd59:
				// Trace: src/VX_popcount.sv:63:70
				sum = 4'd10;
			6'd60:
				// Trace: src/VX_popcount.sv:64:16
				sum = 4'd11;
			6'd61:
				// Trace: src/VX_popcount.sv:64:34
				sum = 4'd12;
			6'd62:
				// Trace: src/VX_popcount.sv:64:52
				sum = 4'd13;
			6'd63:
				// Trace: src/VX_popcount.sv:64:70
				sum = 4'd14;
		endcase
	// Trace: src/VX_popcount.sv:67:5
	assign data_out = sum;
endmodule
module VX_popcount (
	data_in,
	data_out
);
	// Trace: src/VX_popcount.sv:70:15
	parameter MODEL = 1;
	// Trace: src/VX_popcount.sv:71:15
	parameter N = 1;
	// Trace: src/VX_popcount.sv:72:15
	parameter M = $clog2(N + 1);
	// Trace: src/VX_popcount.sv:74:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_popcount.sv:75:5
	output wire [M - 1:0] data_out;
	// Trace: src/VX_popcount.sv:77:5
	function automatic [M - 1:0] sv2v_cast_ABEB2;
		input reg [M - 1:0] inp;
		sv2v_cast_ABEB2 = inp;
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	generate
		if (N == 1) begin : g_passthru
			// Trace: src/VX_popcount.sv:78:9
			assign data_out = data_in;
		end
		else if (N <= 3) begin : g_popcount3
			// Trace: src/VX_popcount.sv:80:9
			reg [2:0] t_in;
			// Trace: src/VX_popcount.sv:81:9
			wire [1:0] t_out;
			// Trace: src/VX_popcount.sv:82:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:83:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:84:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:86:9
			VX_popcount32 pc32(
				.data_in(t_in),
				.data_out(t_out)
			);
			// Trace: src/VX_popcount.sv:87:9
			assign data_out = t_out[M - 1:0];
		end
		else if (N <= 6) begin : g_popcount6
			// Trace: src/VX_popcount.sv:89:9
			reg [5:0] t_in;
			// Trace: src/VX_popcount.sv:90:9
			wire [2:0] t_out;
			// Trace: src/VX_popcount.sv:91:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:92:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:93:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:95:9
			VX_popcount63 pc63(
				.data_in(t_in),
				.data_out(t_out)
			);
			// Trace: src/VX_popcount.sv:96:9
			assign data_out = t_out[M - 1:0];
		end
		else if (N <= 9) begin : g_popcount9
			// Trace: src/VX_popcount.sv:98:9
			reg [8:0] t_in;
			// Trace: src/VX_popcount.sv:99:9
			wire [4:0] t1_out;
			// Trace: src/VX_popcount.sv:100:9
			wire [3:0] t2_out;
			// Trace: src/VX_popcount.sv:101:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:102:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:103:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:105:9
			VX_popcount63 pc63(
				.data_in(t_in[5:0]),
				.data_out(t1_out[2:0])
			);
			// Trace: src/VX_popcount.sv:106:9
			VX_popcount32 pc32(
				.data_in(t_in[8:6]),
				.data_out(t1_out[4:3])
			);
			// Trace: src/VX_popcount.sv:107:9
			VX_sum33 sum33(
				.data_in1(t1_out[2:0]),
				.data_in2({1'b0, t1_out[4:3]}),
				.data_out(t2_out)
			);
			// Trace: src/VX_popcount.sv:108:9
			assign data_out = t2_out[M - 1:0];
		end
		else if (N <= 12) begin : g_popcount12
			// Trace: src/VX_popcount.sv:110:9
			reg [11:0] t_in;
			// Trace: src/VX_popcount.sv:111:9
			wire [5:0] t1_out;
			// Trace: src/VX_popcount.sv:112:9
			wire [3:0] t2_out;
			// Trace: src/VX_popcount.sv:113:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:114:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:115:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:117:9
			VX_popcount63 pc63a(
				.data_in(t_in[5:0]),
				.data_out(t1_out[2:0])
			);
			// Trace: src/VX_popcount.sv:118:9
			VX_popcount63 pc63b(
				.data_in(t_in[11:6]),
				.data_out(t1_out[5:3])
			);
			// Trace: src/VX_popcount.sv:119:9
			VX_sum33 sum33(
				.data_in1(t1_out[2:0]),
				.data_in2(t1_out[5:3]),
				.data_out(t2_out)
			);
			// Trace: src/VX_popcount.sv:120:9
			assign data_out = t2_out[M - 1:0];
		end
		else if (N <= 18) begin : g_popcount18
			// Trace: src/VX_popcount.sv:122:9
			reg [17:0] t_in;
			// Trace: src/VX_popcount.sv:123:9
			wire [8:0] t1_out;
			// Trace: src/VX_popcount.sv:124:9
			wire [5:0] t2_out;
			// Trace: src/VX_popcount.sv:125:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:126:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:127:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:129:9
			VX_popcount63 pc63a(
				.data_in(t_in[5:0]),
				.data_out(t1_out[2:0])
			);
			// Trace: src/VX_popcount.sv:130:9
			VX_popcount63 pc63b(
				.data_in(t_in[11:6]),
				.data_out(t1_out[5:3])
			);
			// Trace: src/VX_popcount.sv:131:9
			VX_popcount63 pc63c(
				.data_in(t_in[17:12]),
				.data_out(t1_out[8:6])
			);
			// Trace: src/VX_popcount.sv:132:9
			VX_popcount32 pc32a(
				.data_in({t1_out[0], t1_out[3], t1_out[6]}),
				.data_out(t2_out[1:0])
			);
			// Trace: src/VX_popcount.sv:133:9
			VX_popcount32 pc32b(
				.data_in({t1_out[1], t1_out[4], t1_out[7]}),
				.data_out(t2_out[3:2])
			);
			// Trace: src/VX_popcount.sv:134:9
			VX_popcount32 pc32c(
				.data_in({t1_out[2], t1_out[5], t1_out[8]}),
				.data_out(t2_out[5:4])
			);
			// Trace: src/VX_popcount.sv:135:9
			assign data_out = ({2'b00, t2_out[1:0]} + {1'b0, t2_out[3:2], 1'b0}) + {t2_out[5:4], 2'b00};
		end
		else if (MODEL == 1) begin : g_model1
			// Trace: src/VX_popcount.sv:137:9
			localparam PN = 1 << $clog2(N);
			// Trace: src/VX_popcount.sv:138:9
			localparam LOGPN = $clog2(PN);
			// Trace: src/VX_popcount.sv:139:9
			wire [M - 1:0] tmp [LOGPN - 1:0][PN - 1:0];
			genvar _gv_j_17;
			for (_gv_j_17 = 0; _gv_j_17 < LOGPN; _gv_j_17 = _gv_j_17 + 1) begin : genblk1
				localparam j = _gv_j_17;
				// Trace: src/VX_popcount.sv:141:13
				localparam D = j + 1;
				// Trace: src/VX_popcount.sv:142:13
				localparam Q = (D < LOGPN ? D + 1 : M);
				genvar _gv_i_166;
				for (_gv_i_166 = 0; _gv_i_166 < (1 << ((LOGPN - j) - 1)); _gv_i_166 = _gv_i_166 + 1) begin : genblk1
					localparam i = _gv_i_166;
					// Trace: src/VX_popcount.sv:144:17
					localparam l = i * 2;
					// Trace: src/VX_popcount.sv:145:17
					localparam r = (i * 2) + 1;
					// Trace: src/VX_popcount.sv:146:17
					wire [Q - 1:0] res;
					if (j == 0) begin : genblk1
						if (r < N) begin : genblk1
							// Trace: src/VX_popcount.sv:149:25
							assign res = data_in[l] + data_in[r];
						end
						else if (l < N) begin : genblk1
							// Trace: src/VX_popcount.sv:151:25
							assign res = sv2v_cast_2(data_in[l]);
						end
						else begin : genblk1
							// Trace: src/VX_popcount.sv:153:25
							assign res = 2'b00;
						end
					end
					else begin : genblk1
						// Trace: src/VX_popcount.sv:156:21
						function automatic [D - 1:0] sv2v_cast_AC9B9;
							input reg [D - 1:0] inp;
							sv2v_cast_AC9B9 = inp;
						endfunction
						assign res = sv2v_cast_AC9B9(tmp[j - 1][l]) + sv2v_cast_AC9B9(tmp[j - 1][r]);
					end
					// Trace: src/VX_popcount.sv:158:17
					assign tmp[j][i] = sv2v_cast_ABEB2(res);
				end
			end
			// Trace: src/VX_popcount.sv:161:9
			assign data_out = tmp[LOGPN - 1][0];
		end
		else begin : g_model2
			// Trace: src/VX_popcount.sv:163:9
			reg [M - 1:0] cnt_w;
			// Trace: src/VX_popcount.sv:164:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:165:13
				cnt_w = 1'sb0;
				// Trace: src/VX_popcount.sv:166:13
				begin : sv2v_autoblock_1
					// Trace: src/VX_popcount.sv:166:18
					integer i;
					// Trace: src/VX_popcount.sv:166:18
					for (i = 0; i < N; i = i + 1)
						begin
							// Trace: src/VX_popcount.sv:167:17
							cnt_w = cnt_w + sv2v_cast_ABEB2(data_in[i]);
						end
				end
			end
			// Trace: src/VX_popcount.sv:170:9
			assign data_out = cnt_w;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_cache_wrap
module VX_elastic_adapter (
	clk,
	reset,
	valid_in,
	ready_in,
	ready_out,
	valid_out,
	busy,
	strobe
);
	// Trace: src/VX_elastic_adapter.sv:2:5
	input wire clk;
	// Trace: src/VX_elastic_adapter.sv:3:5
	input wire reset;
	// Trace: src/VX_elastic_adapter.sv:4:5
	input wire valid_in;
	// Trace: src/VX_elastic_adapter.sv:5:5
	output wire ready_in;
	// Trace: src/VX_elastic_adapter.sv:6:5
	input wire ready_out;
	// Trace: src/VX_elastic_adapter.sv:7:5
	output wire valid_out;
	// Trace: src/VX_elastic_adapter.sv:8:5
	input wire busy;
	// Trace: src/VX_elastic_adapter.sv:9:5
	output wire strobe;
	// Trace: src/VX_elastic_adapter.sv:11:5
	wire push = valid_in && ready_in;
	// Trace: src/VX_elastic_adapter.sv:12:5
	wire pop = valid_out && ready_out;
	// Trace: src/VX_elastic_adapter.sv:13:5
	reg loaded;
	// Trace: src/VX_elastic_adapter.sv:14:5
	always @(posedge clk)
		// Trace: src/VX_elastic_adapter.sv:15:9
		if (reset)
			// Trace: src/VX_elastic_adapter.sv:16:13
			loaded <= 0;
		else begin
			// Trace: src/VX_elastic_adapter.sv:18:13
			if (push)
				// Trace: src/VX_elastic_adapter.sv:19:17
				loaded <= 1;
			if (pop)
				// Trace: src/VX_elastic_adapter.sv:22:17
				loaded <= 0;
		end
	// Trace: src/VX_elastic_adapter.sv:26:5
	assign ready_in = ~loaded;
	// Trace: src/VX_elastic_adapter.sv:27:5
	assign valid_out = loaded && ~busy;
	// Trace: src/VX_elastic_adapter.sv:28:5
	assign strobe = push;
endmodule
module VX_bank_flush (
	clk,
	reset,
	flush_begin,
	flush_end,
	flush_init,
	flush_valid,
	flush_line,
	flush_way,
	flush_ready,
	mshr_empty,
	bank_empty
);
	// Trace: src/VX_bank_flush.sv:2:15
	parameter BANK_ID = 0;
	// Trace: src/VX_bank_flush.sv:3:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_bank_flush.sv:4:15
	parameter LINE_SIZE = 64;
	// Trace: src/VX_bank_flush.sv:5:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_bank_flush.sv:6:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_bank_flush.sv:7:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_bank_flush.sv:9:5
	input wire clk;
	// Trace: src/VX_bank_flush.sv:10:5
	input wire reset;
	// Trace: src/VX_bank_flush.sv:11:5
	input wire flush_begin;
	// Trace: src/VX_bank_flush.sv:12:5
	output wire flush_end;
	// Trace: src/VX_bank_flush.sv:13:5
	output wire flush_init;
	// Trace: src/VX_bank_flush.sv:14:5
	output wire flush_valid;
	// Trace: src/VX_bank_flush.sv:15:5
	output wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] flush_line;
	// Trace: src/VX_bank_flush.sv:16:5
	output wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] flush_way;
	// Trace: src/VX_bank_flush.sv:17:5
	input wire flush_ready;
	// Trace: src/VX_bank_flush.sv:18:5
	input wire mshr_empty;
	// Trace: src/VX_bank_flush.sv:19:5
	input wire bank_empty;
	// Trace: src/VX_bank_flush.sv:21:5
	localparam CTR_WIDTH = $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) + (WRITEBACK ? $clog2(NUM_WAYS) : 0);
	// Trace: src/VX_bank_flush.sv:22:5
	localparam STATE_IDLE = 0;
	// Trace: src/VX_bank_flush.sv:23:5
	localparam STATE_INIT = 1;
	// Trace: src/VX_bank_flush.sv:24:5
	localparam STATE_WAIT1 = 2;
	// Trace: src/VX_bank_flush.sv:25:5
	localparam STATE_FLUSH = 3;
	// Trace: src/VX_bank_flush.sv:26:5
	localparam STATE_WAIT2 = 4;
	// Trace: src/VX_bank_flush.sv:27:5
	localparam STATE_DONE = 5;
	// Trace: src/VX_bank_flush.sv:28:5
	reg [2:0] state;
	reg [2:0] state_n;
	// Trace: src/VX_bank_flush.sv:29:5
	reg [CTR_WIDTH - 1:0] counter;
	// Trace: src/VX_bank_flush.sv:30:5
	always @(*) begin
		// Trace: src/VX_bank_flush.sv:31:9
		state_n = state;
		// Trace: src/VX_bank_flush.sv:32:9
		case (state)
			default:
				// Trace: src/VX_bank_flush.sv:34:17
				if (flush_begin)
					// Trace: src/VX_bank_flush.sv:35:21
					state_n = STATE_WAIT1;
			STATE_INIT:
				// Trace: src/VX_bank_flush.sv:39:17
				if (counter == ((2 ** $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))
					// Trace: src/VX_bank_flush.sv:40:21
					state_n = STATE_IDLE;
			STATE_WAIT1:
				// Trace: src/VX_bank_flush.sv:44:17
				if (mshr_empty)
					// Trace: src/VX_bank_flush.sv:45:21
					state_n = STATE_FLUSH;
			STATE_FLUSH:
				// Trace: src/VX_bank_flush.sv:49:17
				if ((counter == ((2 ** CTR_WIDTH) - 1)) && flush_ready)
					// Trace: src/VX_bank_flush.sv:50:21
					state_n = (BANK_ID == 0 ? STATE_DONE : STATE_WAIT2);
			STATE_WAIT2:
				// Trace: src/VX_bank_flush.sv:54:17
				if (bank_empty)
					// Trace: src/VX_bank_flush.sv:55:21
					state_n = STATE_DONE;
			STATE_DONE:
				// Trace: src/VX_bank_flush.sv:59:17
				state_n = STATE_IDLE;
		endcase
	end
	// Trace: src/VX_bank_flush.sv:63:5
	function automatic signed [CTR_WIDTH - 1:0] sv2v_cast_8E811_signed;
		input reg signed [CTR_WIDTH - 1:0] inp;
		sv2v_cast_8E811_signed = inp;
	endfunction
	always @(posedge clk)
		// Trace: src/VX_bank_flush.sv:64:9
		if (reset) begin
			// Trace: src/VX_bank_flush.sv:65:13
			state <= STATE_INIT;
			// Trace: src/VX_bank_flush.sv:66:13
			counter <= 1'sb0;
		end
		else begin
			// Trace: src/VX_bank_flush.sv:68:13
			state <= state_n;
			// Trace: src/VX_bank_flush.sv:69:13
			if (state != STATE_IDLE) begin
				begin
					// Trace: src/VX_bank_flush.sv:70:17
					if ((state == STATE_INIT) || ((state == STATE_FLUSH) && flush_ready))
						// Trace: src/VX_bank_flush.sv:72:21
						counter <= counter + sv2v_cast_8E811_signed(1);
				end
			end
			else
				// Trace: src/VX_bank_flush.sv:75:17
				counter <= 1'sb0;
		end
	// Trace: src/VX_bank_flush.sv:79:5
	assign flush_end = state == STATE_DONE;
	// Trace: src/VX_bank_flush.sv:80:5
	assign flush_init = state == STATE_INIT;
	// Trace: src/VX_bank_flush.sv:81:5
	assign flush_valid = state == STATE_FLUSH;
	// Trace: src/VX_bank_flush.sv:82:5
	assign flush_line = counter[$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0];
	// Trace: src/VX_bank_flush.sv:83:5
	generate
		if (WRITEBACK && (NUM_WAYS > 1)) begin : g_flush_way
			// Trace: src/VX_bank_flush.sv:84:9
			assign flush_way = counter[$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))+:$clog2(NUM_WAYS)];
		end
		else begin : g_flush_way_all
			// Trace: src/VX_bank_flush.sv:86:9
			assign flush_way = 1'sb0;
		end
	endgenerate
endmodule
module VX_serial_div (
	clk,
	reset,
	strobe,
	busy,
	is_signed,
	numer,
	denom,
	quotient,
	remainder
);
	// Trace: src/VX_serial_div.sv:2:15
	parameter WIDTHN = 32;
	// Trace: src/VX_serial_div.sv:3:15
	parameter WIDTHD = 32;
	// Trace: src/VX_serial_div.sv:4:15
	parameter WIDTHQ = 32;
	// Trace: src/VX_serial_div.sv:5:15
	parameter WIDTHR = 32;
	// Trace: src/VX_serial_div.sv:6:15
	parameter LANES = 1;
	// Trace: src/VX_serial_div.sv:8:5
	input wire clk;
	// Trace: src/VX_serial_div.sv:9:5
	input wire reset;
	// Trace: src/VX_serial_div.sv:10:5
	input wire strobe;
	// Trace: src/VX_serial_div.sv:11:5
	output wire busy;
	// Trace: src/VX_serial_div.sv:12:5
	input wire is_signed;
	// Trace: src/VX_serial_div.sv:13:5
	input wire [(LANES * WIDTHN) - 1:0] numer;
	// Trace: src/VX_serial_div.sv:14:5
	input wire [(LANES * WIDTHD) - 1:0] denom;
	// Trace: src/VX_serial_div.sv:15:5
	output wire [(LANES * WIDTHQ) - 1:0] quotient;
	// Trace: src/VX_serial_div.sv:16:5
	output wire [(LANES * WIDTHR) - 1:0] remainder;
	// Trace: src/VX_serial_div.sv:18:5
	localparam MIN_ND = (WIDTHN < WIDTHD ? WIDTHN : WIDTHD);
	// Trace: src/VX_serial_div.sv:19:5
	localparam CNTRW = $clog2(WIDTHN);
	// Trace: src/VX_serial_div.sv:20:5
	reg [((WIDTHN + MIN_ND) >= 0 ? (LANES * ((WIDTHN + MIN_ND) + 1)) - 1 : (LANES * (1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) - 1)):((WIDTHN + MIN_ND) >= 0 ? 0 : (WIDTHN + MIN_ND) + 0)] working;
	// Trace: src/VX_serial_div.sv:21:5
	reg [(LANES * WIDTHD) - 1:0] denom_r;
	// Trace: src/VX_serial_div.sv:22:5
	wire [(LANES * WIDTHN) - 1:0] numer_qual;
	// Trace: src/VX_serial_div.sv:23:5
	wire [(LANES * WIDTHD) - 1:0] denom_qual;
	// Trace: src/VX_serial_div.sv:24:5
	wire [(WIDTHD >= 0 ? (LANES * (WIDTHD + 1)) - 1 : (LANES * (1 - WIDTHD)) + (WIDTHD - 1)):(WIDTHD >= 0 ? 0 : WIDTHD + 0)] sub_result;
	// Trace: src/VX_serial_div.sv:25:5
	reg [LANES - 1:0] inv_quot;
	reg [LANES - 1:0] inv_rem;
	// Trace: src/VX_serial_div.sv:26:5
	reg [CNTRW - 1:0] cntr;
	// Trace: src/VX_serial_div.sv:27:5
	reg busy_r;
	// Trace: src/VX_serial_div.sv:28:5
	genvar _gv_i_172;
	generate
		for (_gv_i_172 = 0; _gv_i_172 < LANES; _gv_i_172 = _gv_i_172 + 1) begin : g_setup
			localparam i = _gv_i_172;
			// Trace: src/VX_serial_div.sv:29:9
			wire negate_numer = is_signed && numer[(i * WIDTHN) + (WIDTHN - 1)];
			// Trace: src/VX_serial_div.sv:30:9
			wire negate_denom = is_signed && denom[(i * WIDTHD) + (WIDTHD - 1)];
			// Trace: src/VX_serial_div.sv:31:9
			assign numer_qual[i * WIDTHN+:WIDTHN] = (negate_numer ? -$signed(numer[i * WIDTHN+:WIDTHN]) : numer[i * WIDTHN+:WIDTHN]);
			// Trace: src/VX_serial_div.sv:32:9
			assign denom_qual[i * WIDTHD+:WIDTHD] = (negate_denom ? -$signed(denom[i * WIDTHD+:WIDTHD]) : denom[i * WIDTHD+:WIDTHD]);
			// Trace: src/VX_serial_div.sv:33:9
			assign sub_result[(WIDTHD >= 0 ? 0 : WIDTHD) + (i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD))+:(WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)] = working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1))) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1)-:((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)] - denom_r[i * WIDTHD+:WIDTHD];
		end
	endgenerate
	// Trace: src/VX_serial_div.sv:35:5
	function automatic signed [CNTRW - 1:0] sv2v_cast_A86AD_signed;
		input reg signed [CNTRW - 1:0] inp;
		sv2v_cast_A86AD_signed = inp;
	endfunction
	always @(posedge clk) begin
		// Trace: src/VX_serial_div.sv:36:9
		if (reset)
			// Trace: src/VX_serial_div.sv:37:13
			busy_r <= 0;
		else begin
			// Trace: src/VX_serial_div.sv:39:13
			if (strobe)
				// Trace: src/VX_serial_div.sv:40:17
				busy_r <= 1;
			if (busy && (cntr == 0))
				// Trace: src/VX_serial_div.sv:43:17
				busy_r <= 0;
		end
		// Trace: src/VX_serial_div.sv:46:9
		cntr <= cntr - sv2v_cast_A86AD_signed(1);
		if (strobe)
			// Trace: src/VX_serial_div.sv:48:13
			cntr <= sv2v_cast_A86AD_signed(WIDTHN - 1);
	end
	// Trace: src/VX_serial_div.sv:51:5
	genvar _gv_i_173;
	generate
		for (_gv_i_173 = 0; _gv_i_173 < LANES; _gv_i_173 = _gv_i_173 + 1) begin : g_div
			localparam i = _gv_i_173;
			// Trace: src/VX_serial_div.sv:52:9
			always @(posedge clk)
				// Trace: src/VX_serial_div.sv:53:13
				if (strobe) begin
					// Trace: src/VX_serial_div.sv:54:17
					working[((WIDTHN + MIN_ND) >= 0 ? 0 : WIDTHN + MIN_ND) + (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND)))+:((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))] <= {{WIDTHD {1'b0}}, numer_qual[i * WIDTHN+:WIDTHN], 1'b0};
					// Trace: src/VX_serial_div.sv:55:17
					denom_r[i * WIDTHD+:WIDTHD] <= denom_qual[i * WIDTHD+:WIDTHD];
					// Trace: src/VX_serial_div.sv:56:17
					inv_quot[i] <= ((denom[i * WIDTHD+:WIDTHD] != 0) && is_signed) && (numer[(i * WIDTHN) + 31] ^ denom[(i * WIDTHD) + 31]);
					// Trace: src/VX_serial_div.sv:57:17
					inv_rem[i] <= is_signed && numer[(i * WIDTHN) + 31];
				end
				else if (busy_r)
					// Trace: src/VX_serial_div.sv:59:17
					working[((WIDTHN + MIN_ND) >= 0 ? 0 : WIDTHN + MIN_ND) + (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND)))+:((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))] <= (sub_result[(i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)) + (WIDTHD >= 0 ? WIDTHD : WIDTHD - WIDTHD)] ? {working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) - 1 : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) - 1 : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) - 1))) + (WIDTHN + MIN_ND)) - 1)-:WIDTHN + MIN_ND], 1'b0} : {sub_result[(WIDTHD >= 0 ? (i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)) + (WIDTHD >= 0 ? WIDTHD - 1 : WIDTHD - (WIDTHD - 1)) : (((i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)) + (WIDTHD >= 0 ? WIDTHD - 1 : WIDTHD - (WIDTHD - 1))) + WIDTHD) - 1)-:WIDTHD], working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHN - 1 : (WIDTHN + MIN_ND) - (WIDTHN - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHN - 1 : (WIDTHN + MIN_ND) - (WIDTHN - 1))) + WIDTHN) - 1)-:WIDTHN], 1'b1});
		end
	endgenerate
	// Trace: src/VX_serial_div.sv:64:5
	genvar _gv_i_174;
	generate
		for (_gv_i_174 = 0; _gv_i_174 < LANES; _gv_i_174 = _gv_i_174 + 1) begin : g_output
			localparam i = _gv_i_174;
			// Trace: src/VX_serial_div.sv:65:9
			wire [WIDTHQ - 1:0] q = working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHQ - 1 : (WIDTHN + MIN_ND) - (WIDTHQ - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHQ - 1 : (WIDTHN + MIN_ND) - (WIDTHQ - 1))) + WIDTHQ) - 1)-:WIDTHQ];
			// Trace: src/VX_serial_div.sv:66:9
			wire [WIDTHR - 1:0] r = working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1))) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1)-:((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)];
			// Trace: src/VX_serial_div.sv:67:9
			assign quotient[i * WIDTHQ+:WIDTHQ] = (inv_quot[i] ? -$signed(q) : q);
			// Trace: src/VX_serial_div.sv:68:9
			assign remainder[i * WIDTHR+:WIDTHR] = (inv_rem[i] ? -$signed(r) : r);
		end
	endgenerate
	// Trace: src/VX_serial_div.sv:70:5
	assign busy = busy_r;
endmodule
// removed interface: VX_mem_perf_if
// removed module with interface ports: VX_scoreboard
// removed interface: VX_lsu_mem_if
module VX_index_buffer (
	clk,
	reset,
	write_addr,
	write_data,
	acquire_en,
	read_addr,
	read_data,
	release_en,
	empty,
	full
);
	// Trace: src/VX_index_buffer.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_index_buffer.sv:3:15
	parameter SIZE = 1;
	// Trace: src/VX_index_buffer.sv:4:15
	parameter LUTRAM = 0;
	// Trace: src/VX_index_buffer.sv:5:15
	parameter ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
	// Trace: src/VX_index_buffer.sv:7:5
	input wire clk;
	// Trace: src/VX_index_buffer.sv:8:5
	input wire reset;
	// Trace: src/VX_index_buffer.sv:9:5
	output wire [ADDRW - 1:0] write_addr;
	// Trace: src/VX_index_buffer.sv:10:5
	input wire [DATAW - 1:0] write_data;
	// Trace: src/VX_index_buffer.sv:11:5
	input wire acquire_en;
	// Trace: src/VX_index_buffer.sv:12:5
	input wire [ADDRW - 1:0] read_addr;
	// Trace: src/VX_index_buffer.sv:13:5
	output wire [DATAW - 1:0] read_data;
	// Trace: src/VX_index_buffer.sv:14:5
	input wire release_en;
	// Trace: src/VX_index_buffer.sv:15:5
	output wire empty;
	// Trace: src/VX_index_buffer.sv:16:5
	output wire full;
	// Trace: src/VX_index_buffer.sv:18:5
	VX_allocator #(.SIZE(SIZE)) allocator(
		.clk(clk),
		.reset(reset),
		.acquire_en(acquire_en),
		.acquire_addr(write_addr),
		.release_en(release_en),
		.release_addr(read_addr),
		.empty(empty),
		.full(full)
	);
	// Trace: src/VX_index_buffer.sv:30:5
	VX_dp_ram #(
		.DATAW(DATAW),
		.SIZE(SIZE),
		.LUTRAM(LUTRAM),
		.RDW_MODE("W")
	) data_table(
		.clk(clk),
		.reset(reset),
		.read(1'b1),
		.write(acquire_en),
		.wren(1'b1),
		.waddr(write_addr),
		.wdata(write_data),
		.raddr(read_addr),
		.rdata(read_data)
	);
endmodule
module VX_pipe_register (
	clk,
	reset,
	enable,
	data_in,
	data_out
);
	// Trace: src/VX_pipe_register.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_pipe_register.sv:3:15
	parameter RESETW = 0;
	// Trace: src/VX_pipe_register.sv:4:15
	parameter [(RESETW > 0 ? RESETW : 1) - 1:0] INIT_VALUE = {(RESETW > 0 ? RESETW : 1) {1'b0}};
	// Trace: src/VX_pipe_register.sv:5:15
	parameter DEPTH = 1;
	// Trace: src/VX_pipe_register.sv:7:5
	input wire clk;
	// Trace: src/VX_pipe_register.sv:8:5
	input wire reset;
	// Trace: src/VX_pipe_register.sv:9:5
	input wire enable;
	// Trace: src/VX_pipe_register.sv:10:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_pipe_register.sv:11:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_pipe_register.sv:13:5
	generate
		if (DEPTH == 0) begin : g_passthru
			// Trace: src/VX_pipe_register.sv:14:9
			assign data_out = data_in;
		end
		else if (DEPTH == 1) begin : g_depth1
			if (RESETW == 0) begin : g_no_reset
				// Trace: src/VX_pipe_register.sv:17:13
				reg [DATAW - 1:0] value;
				// Trace: src/VX_pipe_register.sv:18:13
				always @(posedge clk)
					// Trace: src/VX_pipe_register.sv:19:17
					if (enable)
						// Trace: src/VX_pipe_register.sv:20:21
						value <= data_in;
				// Trace: src/VX_pipe_register.sv:23:13
				assign data_out = value;
			end
			else if (RESETW < DATAW) begin : g_partial_reset
				// Trace: src/VX_pipe_register.sv:25:13
				reg [(DATAW - RESETW) - 1:0] value_d;
				// Trace: src/VX_pipe_register.sv:26:13
				reg [RESETW - 1:0] value_r;
				// Trace: src/VX_pipe_register.sv:27:13
				always @(posedge clk)
					// Trace: src/VX_pipe_register.sv:28:17
					if (reset)
						// Trace: src/VX_pipe_register.sv:29:21
						value_r <= INIT_VALUE;
					else if (enable)
						// Trace: src/VX_pipe_register.sv:31:21
						value_r <= data_in[DATAW - 1:DATAW - RESETW];
				// Trace: src/VX_pipe_register.sv:34:13
				always @(posedge clk)
					// Trace: src/VX_pipe_register.sv:35:17
					if (enable)
						// Trace: src/VX_pipe_register.sv:36:21
						value_d <= data_in[(DATAW - RESETW) - 1:0];
				// Trace: src/VX_pipe_register.sv:39:13
				assign data_out = {value_r, value_d};
			end
			else begin : g_full_reset
				// Trace: src/VX_pipe_register.sv:41:13
				reg [DATAW - 1:0] value;
				// Trace: src/VX_pipe_register.sv:42:13
				always @(posedge clk)
					// Trace: src/VX_pipe_register.sv:43:17
					if (reset)
						// Trace: src/VX_pipe_register.sv:44:21
						value <= INIT_VALUE;
					else if (enable)
						// Trace: src/VX_pipe_register.sv:46:21
						value <= data_in;
				// Trace: src/VX_pipe_register.sv:49:13
				assign data_out = value;
			end
		end
		else begin : g_recursive
			// Trace: src/VX_pipe_register.sv:52:9
			wire [(DEPTH >= 0 ? ((DEPTH + 1) * DATAW) - 1 : ((1 - DEPTH) * DATAW) + ((DEPTH * DATAW) - 1)):(DEPTH >= 0 ? 0 : DEPTH * DATAW)] data_delayed;
			// Trace: src/VX_pipe_register.sv:53:9
			assign data_delayed[(DEPTH >= 0 ? 0 : DEPTH) * DATAW+:DATAW] = data_in;
			genvar _gv_i_177;
			for (_gv_i_177 = 1; _gv_i_177 <= DEPTH; _gv_i_177 = _gv_i_177 + 1) begin : g_pipe_reg
				localparam i = _gv_i_177;
				// Trace: src/VX_pipe_register.sv:55:13
				VX_pipe_register #(
					.DATAW(DATAW),
					.RESETW(RESETW),
					.INIT_VALUE(INIT_VALUE)
				) pipe_reg(
					.clk(clk),
					.reset(reset),
					.enable(enable),
					.data_in(data_delayed[(DEPTH >= 0 ? i - 1 : DEPTH - (i - 1)) * DATAW+:DATAW]),
					.data_out(data_delayed[(DEPTH >= 0 ? i : DEPTH - i) * DATAW+:DATAW])
				);
			end
			// Trace: src/VX_pipe_register.sv:67:9
			assign data_out = data_delayed[(DEPTH >= 0 ? DEPTH : DEPTH - DEPTH) * DATAW+:DATAW];
		end
	endgenerate
endmodule
// removed module with interface ports: VX_fpu_unit
module VX_cache_bank (
	clk,
	reset,
	core_req_valid,
	core_req_addr,
	core_req_rw,
	core_req_wsel,
	core_req_byteen,
	core_req_data,
	core_req_tag,
	core_req_idx,
	core_req_flags,
	core_req_ready,
	core_rsp_valid,
	core_rsp_data,
	core_rsp_tag,
	core_rsp_idx,
	core_rsp_ready,
	mem_req_valid,
	mem_req_addr,
	mem_req_rw,
	mem_req_byteen,
	mem_req_data,
	mem_req_tag,
	mem_req_flags,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready,
	flush_begin,
	flush_uuid,
	flush_end
);
	// Trace: src/VX_cache_bank.sv:2:16
	parameter INSTANCE_ID = "";
	// Trace: src/VX_cache_bank.sv:3:15
	parameter BANK_ID = 0;
	// Trace: src/VX_cache_bank.sv:4:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_cache_bank.sv:5:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_cache_bank.sv:6:15
	parameter LINE_SIZE = 16;
	// Trace: src/VX_cache_bank.sv:7:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_bank.sv:8:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_bank.sv:9:15
	parameter WORD_SIZE = 4;
	// Trace: src/VX_cache_bank.sv:10:15
	parameter CRSQ_SIZE = 1;
	// Trace: src/VX_cache_bank.sv:11:15
	parameter MSHR_SIZE = 1;
	// Trace: src/VX_cache_bank.sv:12:15
	parameter MREQ_SIZE = 1;
	// Trace: src/VX_cache_bank.sv:13:15
	parameter WRITE_ENABLE = 1;
	// Trace: src/VX_cache_bank.sv:14:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_cache_bank.sv:15:15
	parameter DIRTY_BYTES = 0;
	// Trace: src/VX_cache_bank.sv:16:15
	parameter REPL_POLICY = 1;
	// Trace: src/VX_cache_bank.sv:17:15
	parameter UUID_WIDTH = 0;
	// Trace: src/VX_cache_bank.sv:18:15
	parameter TAG_WIDTH = UUID_WIDTH + 1;
	// Trace: src/VX_cache_bank.sv:19:15
	parameter FLAGS_WIDTH = 0;
	// Trace: src/VX_cache_bank.sv:20:15
	parameter CORE_OUT_REG = 0;
	// Trace: src/VX_cache_bank.sv:21:15
	parameter MEM_OUT_REG = 0;
	// Trace: src/VX_cache_bank.sv:22:15
	parameter MSHR_ADDR_WIDTH = (MSHR_SIZE > 1 ? $clog2(MSHR_SIZE) : 1);
	// Trace: src/VX_cache_bank.sv:23:15
	parameter MEM_TAG_WIDTH = UUID_WIDTH + MSHR_ADDR_WIDTH;
	// Trace: src/VX_cache_bank.sv:24:15
	parameter REQ_SEL_WIDTH = ($clog2(NUM_REQS) > 0 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_cache_bank.sv:25:15
	parameter WORD_SEL_WIDTH = ($clog2(LINE_SIZE / WORD_SIZE) > 0 ? $clog2(LINE_SIZE / WORD_SIZE) : 1);
	// Trace: src/VX_cache_bank.sv:27:5
	input wire clk;
	// Trace: src/VX_cache_bank.sv:28:5
	input wire reset;
	// Trace: src/VX_cache_bank.sv:29:5
	input wire core_req_valid;
	// Trace: src/VX_cache_bank.sv:30:5
	input wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] core_req_addr;
	// Trace: src/VX_cache_bank.sv:31:5
	input wire core_req_rw;
	// Trace: src/VX_cache_bank.sv:32:5
	input wire [WORD_SEL_WIDTH - 1:0] core_req_wsel;
	// Trace: src/VX_cache_bank.sv:33:5
	input wire [WORD_SIZE - 1:0] core_req_byteen;
	// Trace: src/VX_cache_bank.sv:34:5
	input wire [(8 * WORD_SIZE) - 1:0] core_req_data;
	// Trace: src/VX_cache_bank.sv:35:5
	input wire [TAG_WIDTH - 1:0] core_req_tag;
	// Trace: src/VX_cache_bank.sv:36:5
	input wire [REQ_SEL_WIDTH - 1:0] core_req_idx;
	// Trace: src/VX_cache_bank.sv:37:5
	input wire [(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) - 1:0] core_req_flags;
	// Trace: src/VX_cache_bank.sv:38:5
	output wire core_req_ready;
	// Trace: src/VX_cache_bank.sv:39:5
	output wire core_rsp_valid;
	// Trace: src/VX_cache_bank.sv:40:5
	output wire [(8 * WORD_SIZE) - 1:0] core_rsp_data;
	// Trace: src/VX_cache_bank.sv:41:5
	output wire [TAG_WIDTH - 1:0] core_rsp_tag;
	// Trace: src/VX_cache_bank.sv:42:5
	output wire [REQ_SEL_WIDTH - 1:0] core_rsp_idx;
	// Trace: src/VX_cache_bank.sv:43:5
	input wire core_rsp_ready;
	// Trace: src/VX_cache_bank.sv:44:5
	output wire mem_req_valid;
	// Trace: src/VX_cache_bank.sv:45:5
	output wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mem_req_addr;
	// Trace: src/VX_cache_bank.sv:46:5
	output wire mem_req_rw;
	// Trace: src/VX_cache_bank.sv:47:5
	output wire [LINE_SIZE - 1:0] mem_req_byteen;
	// Trace: src/VX_cache_bank.sv:48:5
	output wire [(8 * LINE_SIZE) - 1:0] mem_req_data;
	// Trace: src/VX_cache_bank.sv:49:5
	output wire [MEM_TAG_WIDTH - 1:0] mem_req_tag;
	// Trace: src/VX_cache_bank.sv:50:5
	output wire [(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) - 1:0] mem_req_flags;
	// Trace: src/VX_cache_bank.sv:51:5
	input wire mem_req_ready;
	// Trace: src/VX_cache_bank.sv:52:5
	input wire mem_rsp_valid;
	// Trace: src/VX_cache_bank.sv:53:5
	input wire [(8 * LINE_SIZE) - 1:0] mem_rsp_data;
	// Trace: src/VX_cache_bank.sv:54:5
	input wire [MEM_TAG_WIDTH - 1:0] mem_rsp_tag;
	// Trace: src/VX_cache_bank.sv:55:5
	output wire mem_rsp_ready;
	// Trace: src/VX_cache_bank.sv:56:5
	input wire flush_begin;
	// Trace: src/VX_cache_bank.sv:57:5
	input wire [(UUID_WIDTH > 0 ? UUID_WIDTH : 1) - 1:0] flush_uuid;
	// Trace: src/VX_cache_bank.sv:58:5
	output wire flush_end;
	// Trace: src/VX_cache_bank.sv:60:5
	localparam PIPELINE_STAGES = 2;
	// Trace: src/VX_cache_bank.sv:61:5
	wire [(UUID_WIDTH > 0 ? UUID_WIDTH : 1) - 1:0] req_uuid_sel;
	wire [(UUID_WIDTH > 0 ? UUID_WIDTH : 1) - 1:0] req_uuid_st0;
	wire [(UUID_WIDTH > 0 ? UUID_WIDTH : 1) - 1:0] req_uuid_st1;
	// Trace: src/VX_cache_bank.sv:62:5
	wire crsp_queue_stall;
	// Trace: src/VX_cache_bank.sv:63:5
	wire mshr_alm_full;
	// Trace: src/VX_cache_bank.sv:64:5
	wire mreq_queue_empty;
	// Trace: src/VX_cache_bank.sv:65:5
	wire mreq_queue_alm_full;
	// Trace: src/VX_cache_bank.sv:66:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mem_rsp_addr;
	// Trace: src/VX_cache_bank.sv:67:5
	wire replay_valid;
	// Trace: src/VX_cache_bank.sv:68:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] replay_addr;
	// Trace: src/VX_cache_bank.sv:69:5
	wire replay_rw;
	// Trace: src/VX_cache_bank.sv:70:5
	wire [WORD_SEL_WIDTH - 1:0] replay_wsel;
	// Trace: src/VX_cache_bank.sv:71:5
	wire [WORD_SIZE - 1:0] replay_byteen;
	// Trace: src/VX_cache_bank.sv:72:5
	wire [(8 * WORD_SIZE) - 1:0] replay_data;
	// Trace: src/VX_cache_bank.sv:73:5
	wire [TAG_WIDTH - 1:0] replay_tag;
	// Trace: src/VX_cache_bank.sv:74:5
	wire [REQ_SEL_WIDTH - 1:0] replay_idx;
	// Trace: src/VX_cache_bank.sv:75:5
	wire [MSHR_ADDR_WIDTH - 1:0] replay_id;
	// Trace: src/VX_cache_bank.sv:76:5
	wire replay_ready;
	// Trace: src/VX_cache_bank.sv:77:5
	wire valid_sel;
	wire valid_st0;
	wire valid_st1;
	// Trace: src/VX_cache_bank.sv:78:5
	wire is_init_st0;
	// Trace: src/VX_cache_bank.sv:79:5
	wire is_creq_st0;
	wire is_creq_st1;
	// Trace: src/VX_cache_bank.sv:80:5
	wire is_fill_st0;
	wire is_fill_st1;
	// Trace: src/VX_cache_bank.sv:81:5
	wire is_flush_st0;
	wire is_flush_st1;
	// Trace: src/VX_cache_bank.sv:82:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] flush_way_st0;
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] evict_way_st0;
	// Trace: src/VX_cache_bank.sv:83:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] way_idx_st0;
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] way_idx_st1;
	// Trace: src/VX_cache_bank.sv:84:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_sel;
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_st0;
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_st1;
	// Trace: src/VX_cache_bank.sv:85:5
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx_st0;
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx_st1;
	// Trace: src/VX_cache_bank.sv:86:5
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] line_tag_st0;
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] line_tag_st1;
	// Trace: src/VX_cache_bank.sv:87:5
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] evict_tag_st0;
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] evict_tag_st1;
	// Trace: src/VX_cache_bank.sv:88:5
	wire rw_sel;
	wire rw_st0;
	wire rw_st1;
	// Trace: src/VX_cache_bank.sv:89:5
	wire [WORD_SEL_WIDTH - 1:0] word_idx_sel;
	wire [WORD_SEL_WIDTH - 1:0] word_idx_st0;
	wire [WORD_SEL_WIDTH - 1:0] word_idx_st1;
	// Trace: src/VX_cache_bank.sv:90:5
	wire [WORD_SIZE - 1:0] byteen_sel;
	wire [WORD_SIZE - 1:0] byteen_st0;
	wire [WORD_SIZE - 1:0] byteen_st1;
	// Trace: src/VX_cache_bank.sv:91:5
	wire [REQ_SEL_WIDTH - 1:0] req_idx_sel;
	wire [REQ_SEL_WIDTH - 1:0] req_idx_st0;
	wire [REQ_SEL_WIDTH - 1:0] req_idx_st1;
	// Trace: src/VX_cache_bank.sv:92:5
	wire [TAG_WIDTH - 1:0] tag_sel;
	wire [TAG_WIDTH - 1:0] tag_st0;
	wire [TAG_WIDTH - 1:0] tag_st1;
	// Trace: src/VX_cache_bank.sv:93:5
	wire [(8 * WORD_SIZE) - 1:0] write_word_st0;
	wire [(8 * WORD_SIZE) - 1:0] write_word_st1;
	// Trace: src/VX_cache_bank.sv:94:5
	wire [(8 * LINE_SIZE) - 1:0] data_sel;
	wire [(8 * LINE_SIZE) - 1:0] data_st0;
	wire [(8 * LINE_SIZE) - 1:0] data_st1;
	// Trace: src/VX_cache_bank.sv:95:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_id_st0;
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_id_st1;
	// Trace: src/VX_cache_bank.sv:96:5
	wire [MSHR_ADDR_WIDTH - 1:0] replay_id_st0;
	// Trace: src/VX_cache_bank.sv:97:5
	wire is_dirty_st0;
	wire is_dirty_st1;
	// Trace: src/VX_cache_bank.sv:98:5
	wire is_replay_st0;
	wire is_replay_st1;
	// Trace: src/VX_cache_bank.sv:99:5
	wire is_hit_st0;
	wire is_hit_st1;
	// Trace: src/VX_cache_bank.sv:100:5
	wire [(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) - 1:0] flags_sel;
	wire [(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) - 1:0] flags_st0;
	wire [(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) - 1:0] flags_st1;
	// Trace: src/VX_cache_bank.sv:101:5
	wire mshr_pending_st0;
	wire mshr_pending_st1;
	// Trace: src/VX_cache_bank.sv:102:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_previd_st0;
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_previd_st1;
	// Trace: src/VX_cache_bank.sv:103:5
	wire mshr_empty;
	// Trace: src/VX_cache_bank.sv:104:5
	wire flush_valid;
	// Trace: src/VX_cache_bank.sv:105:5
	wire init_valid;
	// Trace: src/VX_cache_bank.sv:106:5
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] flush_sel;
	// Trace: src/VX_cache_bank.sv:107:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] flush_way;
	// Trace: src/VX_cache_bank.sv:108:5
	wire flush_ready;
	// Trace: src/VX_cache_bank.sv:109:5
	wire no_pending_req = (~valid_st0 && ~valid_st1) && mreq_queue_empty;
	// Trace: src/VX_cache_bank.sv:110:5
	VX_bank_flush #(
		.BANK_ID(BANK_ID),
		.CACHE_SIZE(CACHE_SIZE),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_WAYS(NUM_WAYS),
		.WRITEBACK(WRITEBACK)
	) flush_unit(
		.clk(clk),
		.reset(reset),
		.flush_begin(flush_begin),
		.flush_end(flush_end),
		.flush_init(init_valid),
		.flush_valid(flush_valid),
		.flush_line(flush_sel),
		.flush_way(flush_way),
		.flush_ready(flush_ready),
		.mshr_empty(mshr_empty),
		.bank_empty(no_pending_req)
	);
	// Trace: src/VX_cache_bank.sv:130:5
	wire pipe_stall = crsp_queue_stall;
	// Trace: src/VX_cache_bank.sv:131:5
	wire replay_grant = ~init_valid;
	// Trace: src/VX_cache_bank.sv:132:5
	wire replay_enable = replay_grant && replay_valid;
	// Trace: src/VX_cache_bank.sv:133:5
	wire fill_grant = ~init_valid && ~replay_enable;
	// Trace: src/VX_cache_bank.sv:134:5
	wire fill_enable = fill_grant && mem_rsp_valid;
	// Trace: src/VX_cache_bank.sv:135:5
	wire flush_grant = (~init_valid && ~replay_enable) && ~fill_enable;
	// Trace: src/VX_cache_bank.sv:136:5
	wire flush_enable = flush_grant && flush_valid;
	// Trace: src/VX_cache_bank.sv:137:5
	wire creq_grant = ((~init_valid && ~replay_enable) && ~fill_enable) && ~flush_enable;
	// Trace: src/VX_cache_bank.sv:138:5
	wire creq_enable = creq_grant && core_req_valid;
	// Trace: src/VX_cache_bank.sv:139:5
	assign replay_ready = (replay_grant && ~((!WRITEBACK && replay_rw) && mreq_queue_alm_full)) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:142:5
	assign mem_rsp_ready = (fill_grant && ~(WRITEBACK && mreq_queue_alm_full)) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:145:5
	assign flush_ready = (flush_grant && ~(WRITEBACK && mreq_queue_alm_full)) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:148:5
	assign core_req_ready = ((creq_grant && ~mreq_queue_alm_full) && ~mshr_alm_full) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:152:5
	wire init_fire = init_valid;
	// Trace: src/VX_cache_bank.sv:153:5
	wire replay_fire = replay_valid && replay_ready;
	// Trace: src/VX_cache_bank.sv:154:5
	wire mem_rsp_fire = mem_rsp_valid && mem_rsp_ready;
	// Trace: src/VX_cache_bank.sv:155:5
	wire flush_fire = flush_valid && flush_ready;
	// Trace: src/VX_cache_bank.sv:156:5
	wire core_req_fire = core_req_valid && core_req_ready;
	// Trace: src/VX_cache_bank.sv:157:5
	wire [MSHR_ADDR_WIDTH - 1:0] mem_rsp_id = mem_rsp_tag[MSHR_ADDR_WIDTH - 1:0];
	// Trace: src/VX_cache_bank.sv:158:5
	wire [TAG_WIDTH - 1:0] mem_rsp_tag_s;
	// Trace: src/VX_cache_bank.sv:159:5
	function automatic [(TAG_WIDTH - MEM_TAG_WIDTH) - 1:0] sv2v_cast_E6004;
		input reg [(TAG_WIDTH - MEM_TAG_WIDTH) - 1:0] inp;
		sv2v_cast_E6004 = inp;
	endfunction
	generate
		if (TAG_WIDTH > MEM_TAG_WIDTH) begin : g_mem_rsp_tag_s_pad
			// Trace: src/VX_cache_bank.sv:160:9
			assign mem_rsp_tag_s = {mem_rsp_tag, sv2v_cast_E6004(1'b0)};
		end
		else begin : g_mem_rsp_tag_s_cut
			// Trace: src/VX_cache_bank.sv:162:9
			assign mem_rsp_tag_s = mem_rsp_tag[MEM_TAG_WIDTH - 1-:TAG_WIDTH];
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:164:5
	wire [TAG_WIDTH - 1:0] flush_tag;
	// Trace: src/VX_cache_bank.sv:165:5
	function automatic [(TAG_WIDTH - UUID_WIDTH) - 1:0] sv2v_cast_B8F42;
		input reg [(TAG_WIDTH - UUID_WIDTH) - 1:0] inp;
		sv2v_cast_B8F42 = inp;
	endfunction
	generate
		if (UUID_WIDTH != 0) begin : g_flush_tag_uuid
			// Trace: src/VX_cache_bank.sv:166:9
			assign flush_tag = {flush_uuid, sv2v_cast_B8F42(1'b0)};
		end
		else begin : g_flush_tag_0
			// Trace: src/VX_cache_bank.sv:168:9
			assign flush_tag = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:170:5
	assign valid_sel = (((init_fire || replay_fire) || mem_rsp_fire) || flush_fire) || core_req_fire;
	// Trace: src/VX_cache_bank.sv:171:5
	assign rw_sel = (replay_valid ? replay_rw : core_req_rw);
	// Trace: src/VX_cache_bank.sv:172:5
	assign byteen_sel = (replay_valid ? replay_byteen : core_req_byteen);
	// Trace: src/VX_cache_bank.sv:173:5
	function automatic [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] sv2v_cast_9CD28;
		input reg [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] inp;
		sv2v_cast_9CD28 = inp;
	endfunction
	assign addr_sel = (init_valid | flush_valid ? sv2v_cast_9CD28(flush_sel) : (replay_valid ? replay_addr : (mem_rsp_valid ? mem_rsp_addr : core_req_addr)));
	// Trace: src/VX_cache_bank.sv:175:5
	assign word_idx_sel = (replay_valid ? replay_wsel : core_req_wsel);
	// Trace: src/VX_cache_bank.sv:176:5
	assign req_idx_sel = (replay_valid ? replay_idx : core_req_idx);
	// Trace: src/VX_cache_bank.sv:177:5
	assign tag_sel = (init_valid | flush_valid ? (flush_valid ? flush_tag : {TAG_WIDTH {1'sb0}}) : (replay_valid ? replay_tag : (mem_rsp_valid ? mem_rsp_tag_s : core_req_tag)));
	// Trace: src/VX_cache_bank.sv:179:5
	assign flags_sel = (core_req_valid ? core_req_flags : {(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) {1'sb0}});
	// Trace: src/VX_cache_bank.sv:180:5
	generate
		if (WRITE_ENABLE) begin : g_data_sel
			genvar _gv_i_178;
			for (_gv_i_178 = 0; _gv_i_178 < (8 * LINE_SIZE); _gv_i_178 = _gv_i_178 + 1) begin : g_i
				localparam i = _gv_i_178;
				if (i < (8 * WORD_SIZE)) begin : g_lo
					// Trace: src/VX_cache_bank.sv:183:17
					assign data_sel[i] = (replay_valid ? replay_data[i] : (mem_rsp_valid ? mem_rsp_data[i] : core_req_data[i]));
				end
				else begin : g_hi
					// Trace: src/VX_cache_bank.sv:185:17
					assign data_sel[i] = mem_rsp_data[i];
				end
			end
		end
		else begin : g_data_sel_ro
			// Trace: src/VX_cache_bank.sv:189:9
			assign data_sel = mem_rsp_data;
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:191:5
	generate
		if (UUID_WIDTH != 0) begin : g_req_uuid_sel
			// Trace: src/VX_cache_bank.sv:192:9
			assign req_uuid_sel = tag_sel[TAG_WIDTH - 1-:UUID_WIDTH];
		end
		else begin : g_req_uuid_sel_0
			// Trace: src/VX_cache_bank.sv:194:9
			assign req_uuid_sel = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:196:5
	wire is_init_sel = init_valid;
	// Trace: src/VX_cache_bank.sv:197:5
	wire is_creq_sel = creq_enable || replay_enable;
	// Trace: src/VX_cache_bank.sv:198:5
	wire is_fill_sel = fill_enable;
	// Trace: src/VX_cache_bank.sv:199:5
	wire is_flush_sel = flush_enable;
	// Trace: src/VX_cache_bank.sv:200:5
	wire is_replay_sel = replay_enable;
	// Trace: src/VX_cache_bank.sv:201:5
	VX_pipe_register #(
		.DATAW((((((((((6 + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + ($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1)) + ((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS))) + (8 * LINE_SIZE)) + 1) + WORD_SIZE) + WORD_SEL_WIDTH) + REQ_SEL_WIDTH) + TAG_WIDTH) + MSHR_ADDR_WIDTH),
		.RESETW(1)
	) pipe_reg0(
		.clk(clk),
		.reset(reset),
		.enable(~pipe_stall),
		.data_in({valid_sel, is_init_sel, is_fill_sel, is_flush_sel, is_creq_sel, is_replay_sel, flags_sel, flush_way, addr_sel, data_sel, rw_sel, byteen_sel, word_idx_sel, req_idx_sel, tag_sel, replay_id}),
		.data_out({valid_st0, is_init_st0, is_fill_st0, is_flush_st0, is_creq_st0, is_replay_st0, flags_st0, flush_way_st0, addr_st0, data_st0, rw_st0, byteen_st0, word_idx_st0, req_idx_st0, tag_st0, replay_id_st0})
	);
	// Trace: src/VX_cache_bank.sv:211:5
	generate
		if (UUID_WIDTH != 0) begin : g_req_uuid_st0
			// Trace: src/VX_cache_bank.sv:212:9
			assign req_uuid_st0 = tag_st0[TAG_WIDTH - 1-:UUID_WIDTH];
		end
		else begin : g_req_uuid_st0_0
			// Trace: src/VX_cache_bank.sv:214:9
			assign req_uuid_st0 = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:216:5
	wire is_read_st0 = is_creq_st0 && ~rw_st0;
	// Trace: src/VX_cache_bank.sv:217:5
	wire is_write_st0 = is_creq_st0 && rw_st0;
	// Trace: src/VX_cache_bank.sv:218:5
	wire do_init_st0 = valid_st0 && is_init_st0;
	// Trace: src/VX_cache_bank.sv:219:5
	wire do_flush_st0 = valid_st0 && is_flush_st0;
	// Trace: src/VX_cache_bank.sv:220:5
	wire do_read_st0 = valid_st0 && is_read_st0;
	// Trace: src/VX_cache_bank.sv:221:5
	wire do_write_st0 = valid_st0 && is_write_st0;
	// Trace: src/VX_cache_bank.sv:222:5
	wire do_fill_st0 = valid_st0 && is_fill_st0;
	// Trace: src/VX_cache_bank.sv:223:5
	wire is_read_st1 = is_creq_st1 && ~rw_st1;
	// Trace: src/VX_cache_bank.sv:224:5
	wire is_write_st1 = is_creq_st1 && rw_st1;
	// Trace: src/VX_cache_bank.sv:225:5
	wire do_read_st1 = valid_st1 && is_read_st1;
	// Trace: src/VX_cache_bank.sv:226:5
	wire do_write_st1 = valid_st1 && is_write_st1;
	// Trace: src/VX_cache_bank.sv:227:5
	assign line_idx_st0 = addr_st0[$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0];
	// Trace: src/VX_cache_bank.sv:228:5
	assign line_tag_st0 = addr_st0[((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))];
	// Trace: src/VX_cache_bank.sv:229:5
	assign write_word_st0 = data_st0[(8 * WORD_SIZE) - 1:0];
	// Trace: src/VX_cache_bank.sv:230:5
	wire do_lookup_st0 = do_read_st0 || do_write_st0;
	// Trace: src/VX_cache_bank.sv:231:5
	wire do_lookup_st1 = do_read_st1 || do_write_st1;
	// Trace: src/VX_cache_bank.sv:232:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] victim_way_st0;
	// Trace: src/VX_cache_bank.sv:233:5
	wire [NUM_WAYS - 1:0] tag_matches_st0;
	// Trace: src/VX_cache_bank.sv:234:5
	VX_cache_repl #(
		.CACHE_SIZE(CACHE_SIZE),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_WAYS(NUM_WAYS),
		.REPL_POLICY(REPL_POLICY)
	) cache_repl(
		.clk(clk),
		.reset(reset),
		.stall(pipe_stall),
		.hit_valid((do_lookup_st1 && is_hit_st1) && ~pipe_stall),
		.hit_line(line_idx_st1),
		.hit_way(way_idx_st1),
		.repl_valid(do_fill_st0 && ~pipe_stall),
		.repl_line(line_idx_st0),
		.repl_way(victim_way_st0)
	);
	// Trace: src/VX_cache_bank.sv:251:5
	assign evict_way_st0 = (is_fill_st0 ? victim_way_st0 : flush_way_st0);
	// Trace: src/VX_cache_bank.sv:252:5
	VX_cache_tags #(
		.CACHE_SIZE(CACHE_SIZE),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_WAYS(NUM_WAYS),
		.WORD_SIZE(WORD_SIZE),
		.WRITEBACK(WRITEBACK)
	) cache_tags(
		.clk(clk),
		.reset(reset),
		.init(do_init_st0),
		.flush(do_flush_st0 && ~pipe_stall),
		.fill(do_fill_st0 && ~pipe_stall),
		.read(do_read_st0 && ~pipe_stall),
		.write(do_write_st0 && ~pipe_stall),
		.line_idx(line_idx_st0),
		.line_tag(line_tag_st0),
		.evict_way(evict_way_st0),
		.tag_matches(tag_matches_st0),
		.evict_dirty(is_dirty_st0),
		.evict_tag(evict_tag_st0)
	);
	// Trace: src/VX_cache_bank.sv:274:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] hit_idx_st0;
	// Trace: src/VX_cache_bank.sv:275:5
	VX_onehot_encoder #(.N(NUM_WAYS)) way_idx_enc(
		.data_in(tag_matches_st0),
		.data_out(hit_idx_st0),
		.valid_out()
	);
	// Trace: src/VX_cache_bank.sv:282:5
	assign way_idx_st0 = (is_creq_st0 ? hit_idx_st0 : evict_way_st0);
	// Trace: src/VX_cache_bank.sv:283:5
	assign is_hit_st0 = |tag_matches_st0;
	// Trace: src/VX_cache_bank.sv:284:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_alloc_id_st0;
	// Trace: src/VX_cache_bank.sv:285:5
	assign mshr_id_st0 = (is_replay_st0 ? replay_id_st0 : mshr_alloc_id_st0);
	// Trace: src/VX_cache_bank.sv:286:5
	VX_pipe_register #(
		.DATAW(((((((((((((8 + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + ($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1)) + (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))) + (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) + (8 * LINE_SIZE)) + WORD_SIZE) + WORD_SEL_WIDTH) + REQ_SEL_WIDTH) + TAG_WIDTH) + MSHR_ADDR_WIDTH) + MSHR_ADDR_WIDTH) + 1),
		.RESETW(1)
	) pipe_reg1(
		.clk(clk),
		.reset(reset),
		.enable(~pipe_stall),
		.data_in({valid_st0, is_fill_st0, is_flush_st0, is_creq_st0, is_replay_st0, is_dirty_st0, is_hit_st0, rw_st0, flags_st0, way_idx_st0, evict_tag_st0, line_tag_st0, line_idx_st0, data_st0, byteen_st0, word_idx_st0, req_idx_st0, tag_st0, mshr_id_st0, mshr_previd_st0, mshr_pending_st0}),
		.data_out({valid_st1, is_fill_st1, is_flush_st1, is_creq_st1, is_replay_st1, is_dirty_st1, is_hit_st1, rw_st1, flags_st1, way_idx_st1, evict_tag_st1, line_tag_st1, line_idx_st1, data_st1, byteen_st1, word_idx_st1, req_idx_st1, tag_st1, mshr_id_st1, mshr_previd_st1, mshr_pending_st1})
	);
	// Trace: src/VX_cache_bank.sv:296:5
	generate
		if (UUID_WIDTH != 0) begin : g_req_uuid_st1
			// Trace: src/VX_cache_bank.sv:297:9
			assign req_uuid_st1 = tag_st1[TAG_WIDTH - 1-:UUID_WIDTH];
		end
		else begin : g_req_uuid_st1_0
			// Trace: src/VX_cache_bank.sv:299:9
			assign req_uuid_st1 = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:301:5
	assign addr_st1 = {line_tag_st1, line_idx_st1};
	// Trace: src/VX_cache_bank.sv:302:5
	assign write_word_st1 = data_st1[(8 * WORD_SIZE) - 1:0];
	// Trace: src/VX_cache_bank.sv:303:5
	wire [((LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] read_data_st1;
	// Trace: src/VX_cache_bank.sv:304:5
	wire [LINE_SIZE - 1:0] evict_byteen_st1;
	// Trace: src/VX_cache_bank.sv:305:5
	VX_cache_data #(
		.CACHE_SIZE(CACHE_SIZE),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_WAYS(NUM_WAYS),
		.WORD_SIZE(WORD_SIZE),
		.WRITE_ENABLE(WRITE_ENABLE),
		.WRITEBACK(WRITEBACK),
		.DIRTY_BYTES(DIRTY_BYTES)
	) cache_data(
		.clk(clk),
		.reset(reset),
		.stall(pipe_stall),
		.init(do_init_st0),
		.fill(do_fill_st0 && ~pipe_stall),
		.flush(do_flush_st0 && ~pipe_stall),
		.read(do_read_st0 && ~pipe_stall),
		.write(do_write_st0 && ~pipe_stall),
		.evict_way(evict_way_st0),
		.tag_matches(tag_matches_st0),
		.line_idx(line_idx_st0),
		.fill_data(data_st0),
		.write_word(write_word_st0),
		.word_idx(word_idx_st0),
		.write_byteen(byteen_st0),
		.way_idx_r(way_idx_st1),
		.read_data(read_data_st1),
		.evict_byteen(evict_byteen_st1)
	);
	// Trace: src/VX_cache_bank.sv:334:5
	wire mshr_allocate_st0 = (valid_st0 && is_creq_st0) && ~is_replay_st0;
	// Trace: src/VX_cache_bank.sv:335:5
	wire mshr_finalize_st1 = (valid_st1 && is_creq_st1) && ~is_replay_st1;
	// Trace: src/VX_cache_bank.sv:336:5
	wire mshr_release_st1;
	// Trace: src/VX_cache_bank.sv:337:5
	generate
		if (WRITEBACK) begin : g_mshr_release
			// Trace: src/VX_cache_bank.sv:338:9
			assign mshr_release_st1 = is_hit_st1;
		end
		else begin : g_mshr_release_ro
			// Trace: src/VX_cache_bank.sv:340:9
			assign mshr_release_st1 = is_hit_st1 || (rw_st1 && ~mshr_pending_st1);
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:342:5
	wire mshr_release_fire = (mshr_finalize_st1 && mshr_release_st1) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:343:5
	wire [1:0] mshr_dequeue;
	// Trace: src/VX_cache_bank.sv:344:5
	VX_popcount #(
		.N(2),
		.MODEL(1)
	) __mshr_dequeue__(
		.data_in({replay_fire, mshr_release_fire}),
		.data_out(mshr_dequeue)
	);
	// Trace: src/VX_cache_bank.sv:351:5
	VX_pending_size #(
		.SIZE(MSHR_SIZE),
		.DECRW(2)
	) mshr_pending_size(
		.clk(clk),
		.reset(reset),
		.incr(core_req_fire),
		.decr(mshr_dequeue),
		.empty(mshr_empty),
		.alm_empty(),
		.full(mshr_alm_full),
		.alm_full(),
		.size()
	);
	// Trace: src/VX_cache_bank.sv:365:5
	VX_cache_mshr #(
		.INSTANCE_ID(""),
		.BANK_ID(BANK_ID),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.MSHR_SIZE(MSHR_SIZE),
		.WRITEBACK(WRITEBACK),
		.UUID_WIDTH(UUID_WIDTH),
		.DATA_WIDTH((((WORD_SEL_WIDTH + WORD_SIZE) + (8 * WORD_SIZE)) + TAG_WIDTH) + REQ_SEL_WIDTH)
	) cache_mshr(
		.clk(clk),
		.reset(reset),
		.deq_req_uuid(req_uuid_sel),
		.alc_req_uuid(req_uuid_st0),
		.fin_req_uuid(req_uuid_st1),
		.fill_valid(mem_rsp_fire),
		.fill_id(mem_rsp_id),
		.fill_addr(mem_rsp_addr),
		.dequeue_valid(replay_valid),
		.dequeue_addr(replay_addr),
		.dequeue_rw(replay_rw),
		.dequeue_data({replay_wsel, replay_byteen, replay_data, replay_tag, replay_idx}),
		.dequeue_id(replay_id),
		.dequeue_ready(replay_ready),
		.allocate_valid(mshr_allocate_st0 && ~pipe_stall),
		.allocate_addr(addr_st0),
		.allocate_rw(rw_st0),
		.allocate_data({word_idx_st0, byteen_st0, write_word_st0, tag_st0, req_idx_st0}),
		.allocate_id(mshr_alloc_id_st0),
		.allocate_pending(mshr_pending_st0),
		.allocate_previd(mshr_previd_st0),
		.allocate_ready(),
		.finalize_valid(mshr_finalize_st1 && ~pipe_stall),
		.finalize_is_release(mshr_release_st1),
		.finalize_is_pending(mshr_pending_st1),
		.finalize_id(mshr_id_st1),
		.finalize_previd(mshr_previd_st1)
	);
	// Trace: src/VX_cache_bank.sv:403:5
	wire crsp_queue_valid;
	wire crsp_queue_ready;
	// Trace: src/VX_cache_bank.sv:404:5
	wire [(8 * WORD_SIZE) - 1:0] crsp_queue_data;
	// Trace: src/VX_cache_bank.sv:405:5
	wire [REQ_SEL_WIDTH - 1:0] crsp_queue_idx;
	// Trace: src/VX_cache_bank.sv:406:5
	wire [TAG_WIDTH - 1:0] crsp_queue_tag;
	// Trace: src/VX_cache_bank.sv:407:5
	assign crsp_queue_valid = do_read_st1 && is_hit_st1;
	// Trace: src/VX_cache_bank.sv:408:5
	assign crsp_queue_idx = req_idx_st1;
	// Trace: src/VX_cache_bank.sv:409:5
	assign crsp_queue_data = read_data_st1[word_idx_st1 * (8 * WORD_SIZE)+:8 * WORD_SIZE];
	// Trace: src/VX_cache_bank.sv:410:5
	assign crsp_queue_tag = tag_st1;
	// Trace: src/VX_cache_bank.sv:411:5
	VX_elastic_buffer #(
		.DATAW((TAG_WIDTH + (8 * WORD_SIZE)) + REQ_SEL_WIDTH),
		.SIZE(CRSQ_SIZE),
		.OUT_REG(CORE_OUT_REG)
	) core_rsp_queue(
		.clk(clk),
		.reset(reset),
		.valid_in(crsp_queue_valid),
		.ready_in(crsp_queue_ready),
		.data_in({crsp_queue_tag, crsp_queue_data, crsp_queue_idx}),
		.data_out({core_rsp_tag, core_rsp_data, core_rsp_idx}),
		.valid_out(core_rsp_valid),
		.ready_out(core_rsp_ready)
	);
	// Trace: src/VX_cache_bank.sv:425:5
	assign crsp_queue_stall = crsp_queue_valid && ~crsp_queue_ready;
	// Trace: src/VX_cache_bank.sv:426:5
	wire mreq_queue_push;
	wire mreq_queue_pop;
	// Trace: src/VX_cache_bank.sv:427:5
	wire [(8 * LINE_SIZE) - 1:0] mreq_queue_data;
	// Trace: src/VX_cache_bank.sv:428:5
	wire [LINE_SIZE - 1:0] mreq_queue_byteen;
	// Trace: src/VX_cache_bank.sv:429:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mreq_queue_addr;
	// Trace: src/VX_cache_bank.sv:430:5
	wire [MEM_TAG_WIDTH - 1:0] mreq_queue_tag;
	// Trace: src/VX_cache_bank.sv:431:5
	wire mreq_queue_rw;
	// Trace: src/VX_cache_bank.sv:432:5
	wire [(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) - 1:0] mreq_queue_flags;
	// Trace: src/VX_cache_bank.sv:433:5
	wire is_fill_or_flush_st1 = is_fill_st1 || (is_flush_st1 && WRITEBACK);
	// Trace: src/VX_cache_bank.sv:434:5
	wire do_fill_or_flush_st1 = valid_st1 && is_fill_or_flush_st1;
	// Trace: src/VX_cache_bank.sv:435:5
	wire do_writeback_st1 = do_fill_or_flush_st1 && is_dirty_st1;
	// Trace: src/VX_cache_bank.sv:436:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] evict_addr_st1 = {evict_tag_st1, line_idx_st1};
	// Trace: src/VX_cache_bank.sv:437:5
	generate
		if (WRITE_ENABLE) begin : g_mreq_queue
			if (WRITEBACK) begin : g_wb
				if (DIRTY_BYTES) begin : g_dirty_bytes
					// Trace: src/VX_cache_bank.sv:440:17
					wire has_dirty_bytes = |evict_byteen_st1;
				end
				// Trace: src/VX_cache_bank.sv:442:13
				assign mreq_queue_push = (((do_lookup_st1 && ~is_hit_st1) && ~mshr_pending_st1) || do_writeback_st1) && ~pipe_stall;
				// Trace: src/VX_cache_bank.sv:445:13
				assign mreq_queue_addr = (is_fill_or_flush_st1 ? evict_addr_st1 : addr_st1);
				// Trace: src/VX_cache_bank.sv:446:13
				assign mreq_queue_rw = is_fill_or_flush_st1;
				// Trace: src/VX_cache_bank.sv:447:13
				assign mreq_queue_data = read_data_st1;
				// Trace: src/VX_cache_bank.sv:448:13
				assign mreq_queue_byteen = (is_fill_or_flush_st1 ? evict_byteen_st1 : {LINE_SIZE {1'sb1}});
			end
			else begin : g_wt
				// Trace: src/VX_cache_bank.sv:450:13
				wire [LINE_SIZE - 1:0] line_byteen;
				// Trace: src/VX_cache_bank.sv:451:13
				VX_demux #(
					.DATAW(WORD_SIZE),
					.N(LINE_SIZE / WORD_SIZE)
				) byteen_demux(
					.sel_in(word_idx_st1),
					.data_in(byteen_st1),
					.data_out(line_byteen)
				);
				// Trace: src/VX_cache_bank.sv:459:13
				assign mreq_queue_push = (((do_read_st1 && ~is_hit_st1) && ~mshr_pending_st1) || do_write_st1) && ~pipe_stall;
				// Trace: src/VX_cache_bank.sv:462:13
				assign mreq_queue_addr = addr_st1;
				// Trace: src/VX_cache_bank.sv:463:13
				assign mreq_queue_rw = rw_st1;
				// Trace: src/VX_cache_bank.sv:464:13
				assign mreq_queue_data = {LINE_SIZE / WORD_SIZE {write_word_st1}};
				// Trace: src/VX_cache_bank.sv:465:13
				assign mreq_queue_byteen = (rw_st1 ? line_byteen : {LINE_SIZE {1'sb1}});
			end
		end
		else begin : g_mreq_queue_ro
			// Trace: src/VX_cache_bank.sv:468:9
			assign mreq_queue_push = ((do_read_st1 && ~is_hit_st1) && ~mshr_pending_st1) && ~pipe_stall;
			// Trace: src/VX_cache_bank.sv:470:9
			assign mreq_queue_addr = addr_st1;
			// Trace: src/VX_cache_bank.sv:471:9
			assign mreq_queue_rw = 0;
			// Trace: src/VX_cache_bank.sv:472:9
			assign mreq_queue_data = 1'sb0;
			// Trace: src/VX_cache_bank.sv:473:9
			assign mreq_queue_byteen = 1'sb1;
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:475:5
	generate
		if (UUID_WIDTH != 0) begin : g_mreq_queue_tag_uuid
			// Trace: src/VX_cache_bank.sv:476:9
			assign mreq_queue_tag = {req_uuid_st1, mshr_id_st1};
		end
		else begin : g_mreq_queue_tag
			// Trace: src/VX_cache_bank.sv:478:9
			assign mreq_queue_tag = mshr_id_st1;
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:480:5
	assign mreq_queue_pop = mem_req_valid && mem_req_ready;
	// Trace: src/VX_cache_bank.sv:481:5
	assign mreq_queue_flags = flags_st1;
	// Trace: src/VX_cache_bank.sv:482:5
	VX_fifo_queue #(
		.DATAW(((((1 + ((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS))) + LINE_SIZE) + (8 * LINE_SIZE)) + MEM_TAG_WIDTH) + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)),
		.DEPTH(MREQ_SIZE),
		.ALM_FULL(MREQ_SIZE - PIPELINE_STAGES),
		.OUT_REG(MEM_OUT_REG)
	) mem_req_queue(
		.clk(clk),
		.reset(reset),
		.push(mreq_queue_push),
		.pop(mreq_queue_pop),
		.data_in({mreq_queue_rw, mreq_queue_addr, mreq_queue_byteen, mreq_queue_data, mreq_queue_tag, mreq_queue_flags}),
		.data_out({mem_req_rw, mem_req_addr, mem_req_byteen, mem_req_data, mem_req_tag, mem_req_flags}),
		.empty(mreq_queue_empty),
		.alm_full(mreq_queue_alm_full),
		.full(),
		.alm_empty(),
		.size()
	);
	// Trace: src/VX_cache_bank.sv:500:5
	assign mem_req_valid = ~mreq_queue_empty;
endmodule
// removed module with interface ports: VX_cache_bypass
// removed package "VX_fpu_pkg"
module VX_transpose (
	data_in,
	data_out
);
	// Trace: src/VX_transpose.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_transpose.sv:3:15
	parameter N = 1;
	// Trace: src/VX_transpose.sv:4:15
	parameter M = 1;
	// Trace: src/VX_transpose.sv:6:5
	input wire [((N * M) * DATAW) - 1:0] data_in;
	// Trace: src/VX_transpose.sv:7:5
	output wire [((M * N) * DATAW) - 1:0] data_out;
	// Trace: src/VX_transpose.sv:9:5
	genvar _gv_i_183;
	generate
		for (_gv_i_183 = 0; _gv_i_183 < N; _gv_i_183 = _gv_i_183 + 1) begin : g_i
			localparam i = _gv_i_183;
			genvar _gv_j_18;
			for (_gv_j_18 = 0; _gv_j_18 < M; _gv_j_18 = _gv_j_18 + 1) begin : g_j
				localparam j = _gv_j_18;
				// Trace: src/VX_transpose.sv:11:13
				assign data_out[((j * N) + i) * DATAW+:DATAW] = data_in[((i * M) + j) * DATAW+:DATAW];
			end
		end
	endgenerate
endmodule
module VX_stream_switch (
	clk,
	reset,
	sel_in,
	valid_in,
	data_in,
	ready_in,
	valid_out,
	data_out,
	ready_out
);
	// Trace: src/VX_stream_switch.sv:2:15
	parameter NUM_INPUTS = 1;
	// Trace: src/VX_stream_switch.sv:3:15
	parameter NUM_OUTPUTS = 1;
	// Trace: src/VX_stream_switch.sv:4:15
	parameter DATAW = 1;
	// Trace: src/VX_stream_switch.sv:5:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_switch.sv:6:15
	parameter NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
	// Trace: src/VX_stream_switch.sv:7:15
	parameter SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
	// Trace: src/VX_stream_switch.sv:8:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: src/VX_stream_switch.sv:10:5
	input wire clk;
	// Trace: src/VX_stream_switch.sv:11:5
	input wire reset;
	// Trace: src/VX_stream_switch.sv:12:5
	input wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] sel_in;
	// Trace: src/VX_stream_switch.sv:13:5
	input wire [NUM_INPUTS - 1:0] valid_in;
	// Trace: src/VX_stream_switch.sv:14:5
	input wire [(NUM_INPUTS * DATAW) - 1:0] data_in;
	// Trace: src/VX_stream_switch.sv:15:5
	output wire [NUM_INPUTS - 1:0] ready_in;
	// Trace: src/VX_stream_switch.sv:16:5
	output wire [NUM_OUTPUTS - 1:0] valid_out;
	// Trace: src/VX_stream_switch.sv:17:5
	output wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out;
	// Trace: src/VX_stream_switch.sv:18:5
	input wire [NUM_OUTPUTS - 1:0] ready_out;
	// Trace: src/VX_stream_switch.sv:20:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_INPUTS > NUM_OUTPUTS) begin : g_input_select
			genvar _gv_o_9;
			for (_gv_o_9 = 0; _gv_o_9 < NUM_OUTPUTS; _gv_o_9 = _gv_o_9 + 1) begin : g_out_buf
				localparam o = _gv_o_9;
				// Trace: src/VX_stream_switch.sv:22:13
				wire [NUM_REQS - 1:0] valid_in_w;
				// Trace: src/VX_stream_switch.sv:23:13
				wire [(NUM_REQS * DATAW) - 1:0] data_in_w;
				// Trace: src/VX_stream_switch.sv:24:13
				wire [NUM_REQS - 1:0] ready_in_w;
				genvar _gv_r_11;
				for (_gv_r_11 = 0; _gv_r_11 < NUM_REQS; _gv_r_11 = _gv_r_11 + 1) begin : g_r
					localparam r = _gv_r_11;
					// Trace: src/VX_stream_switch.sv:26:17
					localparam i = (r * NUM_OUTPUTS) + o;
					if (i < NUM_INPUTS) begin : g_valid
						// Trace: src/VX_stream_switch.sv:28:21
						assign valid_in_w[r] = valid_in[i];
						// Trace: src/VX_stream_switch.sv:29:21
						assign data_in_w[r * DATAW+:DATAW] = data_in[i * DATAW+:DATAW];
						// Trace: src/VX_stream_switch.sv:30:21
						assign ready_in[i] = ready_in_w[r];
					end
					else begin : g_padding
						// Trace: src/VX_stream_switch.sv:32:21
						assign valid_in_w[r] = 0;
						// Trace: src/VX_stream_switch.sv:33:21
						assign data_in_w[r * DATAW+:DATAW] = 1'sb0;
					end
				end
				// Trace: src/VX_stream_switch.sv:36:13
				VX_elastic_buffer #(
					.DATAW(DATAW),
					.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
					.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
				) out_buf(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_in_w[sel_in[o * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)]]),
					.ready_in(ready_in_w[sel_in[o * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)]]),
					.data_in(data_in_w[sel_in[o * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)] * DATAW+:DATAW]),
					.data_out(data_out[o * DATAW+:DATAW]),
					.valid_out(valid_out[o]),
					.ready_out(ready_out[o])
				);
			end
		end
		else if (NUM_OUTPUTS > NUM_INPUTS) begin : g_output_select
			genvar _gv_i_184;
			for (_gv_i_184 = 0; _gv_i_184 < NUM_INPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_out_buf
				localparam i = _gv_i_184;
				// Trace: src/VX_stream_switch.sv:53:13
				wire [NUM_REQS - 1:0] ready_out_w;
				genvar _gv_r_12;
				for (_gv_r_12 = 0; _gv_r_12 < NUM_REQS; _gv_r_12 = _gv_r_12 + 1) begin : g_r
					localparam r = _gv_r_12;
					// Trace: src/VX_stream_switch.sv:55:17
					localparam o = (r * NUM_INPUTS) + i;
					if (o < NUM_OUTPUTS) begin : g_valid
						// Trace: src/VX_stream_switch.sv:57:21
						wire valid_out_w = valid_in[i] && (sel_in[i * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)] == sv2v_cast_76B5F_signed(r));
						// Trace: src/VX_stream_switch.sv:58:21
						VX_elastic_buffer #(
							.DATAW(DATAW),
							.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
							.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
						) out_buf(
							.clk(clk),
							.reset(reset),
							.valid_in(valid_out_w),
							.ready_in(ready_out_w[r]),
							.data_in(data_in[i * DATAW+:DATAW]),
							.data_out(data_out[o * DATAW+:DATAW]),
							.valid_out(valid_out[o]),
							.ready_out(ready_out[o])
						);
					end
					else begin : g_padding
						// Trace: src/VX_stream_switch.sv:73:21
						assign ready_out_w[r] = 1'sb0;
					end
				end
				// Trace: src/VX_stream_switch.sv:76:13
				assign ready_in[i] = ready_out_w[sel_in[i * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)]];
			end
		end
		else begin : g_passthru
			genvar _gv_i_185;
			for (_gv_i_185 = 0; _gv_i_185 < NUM_OUTPUTS; _gv_i_185 = _gv_i_185 + 1) begin : g_out_buf
				localparam i = _gv_i_185;
				// Trace: src/VX_stream_switch.sv:80:13
				VX_elastic_buffer #(
					.DATAW(DATAW),
					.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
					.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
				) out_buf(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_in[i]),
					.ready_in(ready_in[i]),
					.data_in(data_in[i * DATAW+:DATAW]),
					.data_out(data_out[i * DATAW+:DATAW]),
					.valid_out(valid_out[i]),
					.ready_out(ready_out[i])
				);
			end
		end
	endgenerate
endmodule
// removed module with interface ports: VX_alu_muldiv
module VX_dp_ram (
	clk,
	reset,
	read,
	write,
	wren,
	waddr,
	wdata,
	raddr,
	rdata
);
	// Trace: src/VX_dp_ram.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_dp_ram.sv:3:15
	parameter SIZE = 1;
	// Trace: src/VX_dp_ram.sv:4:15
	parameter WRENW = 1;
	// Trace: src/VX_dp_ram.sv:5:15
	parameter OUT_REG = 0;
	// Trace: src/VX_dp_ram.sv:6:15
	parameter LUTRAM = 0;
	// Trace: src/VX_dp_ram.sv:7:15
	parameter RDW_MODE = "W";
	// Trace: src/VX_dp_ram.sv:8:15
	parameter RADDR_REG = 0;
	// Trace: src/VX_dp_ram.sv:9:15
	parameter RDW_ASSERT = 0;
	// Trace: src/VX_dp_ram.sv:10:15
	parameter RESET_RAM = 0;
	// Trace: src/VX_dp_ram.sv:11:15
	parameter INIT_ENABLE = 0;
	// Trace: src/VX_dp_ram.sv:12:15
	parameter INIT_FILE = "";
	// Trace: src/VX_dp_ram.sv:13:15
	parameter [DATAW - 1:0] INIT_VALUE = 0;
	// Trace: src/VX_dp_ram.sv:14:15
	parameter ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
	// Trace: src/VX_dp_ram.sv:16:5
	input wire clk;
	// Trace: src/VX_dp_ram.sv:17:5
	input wire reset;
	// Trace: src/VX_dp_ram.sv:18:5
	input wire read;
	// Trace: src/VX_dp_ram.sv:19:5
	input wire write;
	// Trace: src/VX_dp_ram.sv:20:5
	input wire [WRENW - 1:0] wren;
	// Trace: src/VX_dp_ram.sv:21:5
	input wire [ADDRW - 1:0] waddr;
	// Trace: src/VX_dp_ram.sv:22:5
	input wire [DATAW - 1:0] wdata;
	// Trace: src/VX_dp_ram.sv:23:5
	input wire [ADDRW - 1:0] raddr;
	// Trace: src/VX_dp_ram.sv:24:5
	output wire [DATAW - 1:0] rdata;
	// Trace: src/VX_dp_ram.sv:26:5
	localparam WSELW = DATAW / WRENW;
	// Trace: src/VX_dp_ram.sv:27:5
	localparam FORCE_BRAM = !LUTRAM && ((SIZE * DATAW) >= 1024);
	// Trace: src/VX_dp_ram.sv:28:5
	generate
		if (OUT_REG) begin : g_sync
			if (FORCE_BRAM) begin : g_bram
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:32:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:35:13
								initial begin
									// Trace: src/VX_dp_ram.sv:35:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:37:13
								initial begin
									// Trace: src/VX_dp_ram.sv:38:17
									begin : sv2v_autoblock_1
										// Trace: src/VX_dp_ram.sv:38:22
										integer i;
										// Trace: src/VX_dp_ram.sv:38:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:39:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:44:21
						reg [ADDRW - 1:0] raddr_r;
						// Trace: src/VX_dp_ram.sv:45:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:46:25
							if (read || write) begin
								// Trace: src/VX_dp_ram.sv:47:29
								if (write)
									// Trace: src/VX_dp_ram.sv:48:33
									begin : sv2v_autoblock_2
										// Trace: src/VX_dp_ram.sv:48:38
										integer i;
										// Trace: src/VX_dp_ram.sv:48:38
										for (i = 0; i < WRENW; i = i + 1)
											begin
												// Trace: src/VX_dp_ram.sv:49:33
												if (wren[i])
													// Trace: src/VX_dp_ram.sv:50:37
													ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
											end
									end
								// Trace: src/VX_dp_ram.sv:54:29
								raddr_r <= raddr;
							end
						// Trace: src/VX_dp_ram.sv:57:21
						assign rdata = ram[raddr_r];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:59:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:62:13
								initial begin
									// Trace: src/VX_dp_ram.sv:62:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:64:13
								initial begin
									// Trace: src/VX_dp_ram.sv:65:17
									begin : sv2v_autoblock_3
										// Trace: src/VX_dp_ram.sv:65:22
										integer i;
										// Trace: src/VX_dp_ram.sv:65:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:66:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:71:21
						reg [ADDRW - 1:0] raddr_r;
						// Trace: src/VX_dp_ram.sv:72:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:73:25
							if (read || write) begin
								// Trace: src/VX_dp_ram.sv:74:29
								if (write)
									// Trace: src/VX_dp_ram.sv:75:33
									ram[waddr] <= wdata;
								// Trace: src/VX_dp_ram.sv:77:29
								raddr_r <= raddr;
							end
						// Trace: src/VX_dp_ram.sv:80:21
						assign rdata = ram[raddr_r];
					end
				end
				else if (RDW_MODE == "R") begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:84:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:87:13
								initial begin
									// Trace: src/VX_dp_ram.sv:87:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:89:13
								initial begin
									// Trace: src/VX_dp_ram.sv:90:17
									begin : sv2v_autoblock_4
										// Trace: src/VX_dp_ram.sv:90:22
										integer i;
										// Trace: src/VX_dp_ram.sv:90:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:91:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:96:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:97:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:98:25
							if (read || write) begin
								// Trace: src/VX_dp_ram.sv:99:29
								if (write)
									// Trace: src/VX_dp_ram.sv:100:33
									begin : sv2v_autoblock_5
										// Trace: src/VX_dp_ram.sv:100:38
										integer i;
										// Trace: src/VX_dp_ram.sv:100:38
										for (i = 0; i < WRENW; i = i + 1)
											begin
												// Trace: src/VX_dp_ram.sv:101:33
												if (wren[i])
													// Trace: src/VX_dp_ram.sv:102:37
													ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
											end
									end
								// Trace: src/VX_dp_ram.sv:106:29
								rdata_r <= ram[raddr];
							end
						// Trace: src/VX_dp_ram.sv:109:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:111:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:114:13
								initial begin
									// Trace: src/VX_dp_ram.sv:114:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:116:13
								initial begin
									// Trace: src/VX_dp_ram.sv:117:17
									begin : sv2v_autoblock_6
										// Trace: src/VX_dp_ram.sv:117:22
										integer i;
										// Trace: src/VX_dp_ram.sv:117:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:118:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:123:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:124:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:125:25
							if (read || write) begin
								// Trace: src/VX_dp_ram.sv:126:29
								if (write)
									// Trace: src/VX_dp_ram.sv:127:33
									ram[waddr] <= wdata;
								// Trace: src/VX_dp_ram.sv:129:29
								rdata_r <= ram[raddr];
							end
						// Trace: src/VX_dp_ram.sv:132:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "U") begin : g_undefined
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:136:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:139:13
								initial begin
									// Trace: src/VX_dp_ram.sv:139:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:141:13
								initial begin
									// Trace: src/VX_dp_ram.sv:142:17
									begin : sv2v_autoblock_7
										// Trace: src/VX_dp_ram.sv:142:22
										integer i;
										// Trace: src/VX_dp_ram.sv:142:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:143:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:148:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:149:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:150:25
							if (write)
								// Trace: src/VX_dp_ram.sv:151:29
								begin : sv2v_autoblock_8
									// Trace: src/VX_dp_ram.sv:151:34
									integer i;
									// Trace: src/VX_dp_ram.sv:151:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:152:33
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:153:37
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_dp_ram.sv:158:29
								rdata_r <= ram[raddr];
						end
						// Trace: src/VX_dp_ram.sv:161:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:163:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:166:13
								initial begin
									// Trace: src/VX_dp_ram.sv:166:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:168:13
								initial begin
									// Trace: src/VX_dp_ram.sv:169:17
									begin : sv2v_autoblock_9
										// Trace: src/VX_dp_ram.sv:169:22
										integer i;
										// Trace: src/VX_dp_ram.sv:169:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:170:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:175:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:176:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:177:25
							if (write)
								// Trace: src/VX_dp_ram.sv:178:29
								ram[waddr] <= wdata;
							if (read)
								// Trace: src/VX_dp_ram.sv:181:29
								rdata_r <= ram[raddr];
						end
						// Trace: src/VX_dp_ram.sv:184:21
						assign rdata = rdata_r;
					end
				end
			end
			else begin : g_auto
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:190:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:193:13
								initial begin
									// Trace: src/VX_dp_ram.sv:193:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:195:13
								initial begin
									// Trace: src/VX_dp_ram.sv:196:17
									begin : sv2v_autoblock_10
										// Trace: src/VX_dp_ram.sv:196:22
										integer i;
										// Trace: src/VX_dp_ram.sv:196:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:197:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:202:21
						reg [ADDRW - 1:0] raddr_r;
						// Trace: src/VX_dp_ram.sv:203:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:204:25
							if (read || write) begin
								// Trace: src/VX_dp_ram.sv:205:29
								if (write)
									// Trace: src/VX_dp_ram.sv:206:33
									begin : sv2v_autoblock_11
										// Trace: src/VX_dp_ram.sv:206:38
										integer i;
										// Trace: src/VX_dp_ram.sv:206:38
										for (i = 0; i < WRENW; i = i + 1)
											begin
												// Trace: src/VX_dp_ram.sv:207:33
												if (wren[i])
													// Trace: src/VX_dp_ram.sv:208:37
													ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
											end
									end
								// Trace: src/VX_dp_ram.sv:212:29
								raddr_r <= raddr;
							end
						// Trace: src/VX_dp_ram.sv:215:21
						assign rdata = ram[raddr_r];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:217:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:220:13
								initial begin
									// Trace: src/VX_dp_ram.sv:220:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:222:13
								initial begin
									// Trace: src/VX_dp_ram.sv:223:17
									begin : sv2v_autoblock_12
										// Trace: src/VX_dp_ram.sv:223:22
										integer i;
										// Trace: src/VX_dp_ram.sv:223:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:224:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:229:21
						reg [ADDRW - 1:0] raddr_r;
						// Trace: src/VX_dp_ram.sv:230:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:231:25
							if (read || write) begin
								// Trace: src/VX_dp_ram.sv:232:29
								if (write)
									// Trace: src/VX_dp_ram.sv:233:33
									ram[waddr] <= wdata;
								// Trace: src/VX_dp_ram.sv:235:29
								raddr_r <= raddr;
							end
						// Trace: src/VX_dp_ram.sv:238:21
						assign rdata = ram[raddr_r];
					end
				end
				else if (RDW_MODE == "R") begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:242:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:245:13
								initial begin
									// Trace: src/VX_dp_ram.sv:245:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:247:13
								initial begin
									// Trace: src/VX_dp_ram.sv:248:17
									begin : sv2v_autoblock_13
										// Trace: src/VX_dp_ram.sv:248:22
										integer i;
										// Trace: src/VX_dp_ram.sv:248:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:249:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:254:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:255:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:256:25
							if (read || write) begin
								// Trace: src/VX_dp_ram.sv:257:29
								if (write)
									// Trace: src/VX_dp_ram.sv:258:33
									begin : sv2v_autoblock_14
										// Trace: src/VX_dp_ram.sv:258:38
										integer i;
										// Trace: src/VX_dp_ram.sv:258:38
										for (i = 0; i < WRENW; i = i + 1)
											begin
												// Trace: src/VX_dp_ram.sv:259:33
												if (wren[i])
													// Trace: src/VX_dp_ram.sv:260:37
													ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
											end
									end
								// Trace: src/VX_dp_ram.sv:264:29
								rdata_r <= ram[raddr];
							end
						// Trace: src/VX_dp_ram.sv:267:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:269:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:272:13
								initial begin
									// Trace: src/VX_dp_ram.sv:272:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:274:13
								initial begin
									// Trace: src/VX_dp_ram.sv:275:17
									begin : sv2v_autoblock_15
										// Trace: src/VX_dp_ram.sv:275:22
										integer i;
										// Trace: src/VX_dp_ram.sv:275:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:276:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:281:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:282:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:283:25
							if (read || write) begin
								// Trace: src/VX_dp_ram.sv:284:29
								if (write)
									// Trace: src/VX_dp_ram.sv:285:33
									ram[waddr] <= wdata;
								// Trace: src/VX_dp_ram.sv:287:29
								rdata_r <= ram[raddr];
							end
						// Trace: src/VX_dp_ram.sv:290:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "U") begin : g_undefined
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:294:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:297:13
								initial begin
									// Trace: src/VX_dp_ram.sv:297:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:299:13
								initial begin
									// Trace: src/VX_dp_ram.sv:300:17
									begin : sv2v_autoblock_16
										// Trace: src/VX_dp_ram.sv:300:22
										integer i;
										// Trace: src/VX_dp_ram.sv:300:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:301:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:306:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:307:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:308:25
							if (write)
								// Trace: src/VX_dp_ram.sv:309:29
								begin : sv2v_autoblock_17
									// Trace: src/VX_dp_ram.sv:309:34
									integer i;
									// Trace: src/VX_dp_ram.sv:309:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:310:33
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:311:37
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_dp_ram.sv:316:29
								rdata_r <= ram[raddr];
						end
						// Trace: src/VX_dp_ram.sv:319:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:321:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:324:13
								initial begin
									// Trace: src/VX_dp_ram.sv:324:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:326:13
								initial begin
									// Trace: src/VX_dp_ram.sv:327:17
									begin : sv2v_autoblock_18
										// Trace: src/VX_dp_ram.sv:327:22
										integer i;
										// Trace: src/VX_dp_ram.sv:327:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:328:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:333:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:334:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:335:25
							if (write)
								// Trace: src/VX_dp_ram.sv:336:29
								ram[waddr] <= wdata;
							if (read)
								// Trace: src/VX_dp_ram.sv:339:29
								rdata_r <= ram[raddr];
						end
						// Trace: src/VX_dp_ram.sv:342:21
						assign rdata = rdata_r;
					end
				end
			end
		end
		else begin : g_async
			if (FORCE_BRAM) begin : g_bram
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:350:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:353:13
								initial begin
									// Trace: src/VX_dp_ram.sv:353:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:355:13
								initial begin
									// Trace: src/VX_dp_ram.sv:356:17
									begin : sv2v_autoblock_19
										// Trace: src/VX_dp_ram.sv:356:22
										integer i;
										// Trace: src/VX_dp_ram.sv:356:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:357:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:362:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:363:25
							if (write)
								// Trace: src/VX_dp_ram.sv:364:29
								begin : sv2v_autoblock_20
									// Trace: src/VX_dp_ram.sv:364:34
									integer i;
									// Trace: src/VX_dp_ram.sv:364:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:365:33
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:366:37
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_dp_ram.sv:371:21
						assign rdata = ram[raddr];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:373:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:376:13
								initial begin
									// Trace: src/VX_dp_ram.sv:376:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:378:13
								initial begin
									// Trace: src/VX_dp_ram.sv:379:17
									begin : sv2v_autoblock_21
										// Trace: src/VX_dp_ram.sv:379:22
										integer i;
										// Trace: src/VX_dp_ram.sv:379:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:380:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:385:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:386:25
							if (write)
								// Trace: src/VX_dp_ram.sv:387:29
								ram[waddr] <= wdata;
						// Trace: src/VX_dp_ram.sv:390:21
						assign rdata = ram[raddr];
					end
				end
				else begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:394:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:397:13
								initial begin
									// Trace: src/VX_dp_ram.sv:397:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:399:13
								initial begin
									// Trace: src/VX_dp_ram.sv:400:17
									begin : sv2v_autoblock_22
										// Trace: src/VX_dp_ram.sv:400:22
										integer i;
										// Trace: src/VX_dp_ram.sv:400:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:401:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:406:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:407:25
							if (write)
								// Trace: src/VX_dp_ram.sv:408:29
								begin : sv2v_autoblock_23
									// Trace: src/VX_dp_ram.sv:408:34
									integer i;
									// Trace: src/VX_dp_ram.sv:408:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:409:33
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:410:37
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_dp_ram.sv:415:21
						assign rdata = ram[raddr];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:417:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:420:13
								initial begin
									// Trace: src/VX_dp_ram.sv:420:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:422:13
								initial begin
									// Trace: src/VX_dp_ram.sv:423:17
									begin : sv2v_autoblock_24
										// Trace: src/VX_dp_ram.sv:423:22
										integer i;
										// Trace: src/VX_dp_ram.sv:423:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:424:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:429:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:430:25
							if (write)
								// Trace: src/VX_dp_ram.sv:431:29
								ram[waddr] <= wdata;
						// Trace: src/VX_dp_ram.sv:434:21
						assign rdata = ram[raddr];
					end
				end
			end
			else begin : g_auto
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:440:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:443:13
								initial begin
									// Trace: src/VX_dp_ram.sv:443:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:445:13
								initial begin
									// Trace: src/VX_dp_ram.sv:446:17
									begin : sv2v_autoblock_25
										// Trace: src/VX_dp_ram.sv:446:22
										integer i;
										// Trace: src/VX_dp_ram.sv:446:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:447:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:452:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:453:25
							if (write)
								// Trace: src/VX_dp_ram.sv:454:29
								begin : sv2v_autoblock_26
									// Trace: src/VX_dp_ram.sv:454:34
									integer i;
									// Trace: src/VX_dp_ram.sv:454:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:455:33
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:456:37
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_dp_ram.sv:461:21
						assign rdata = ram[raddr];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:463:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:466:13
								initial begin
									// Trace: src/VX_dp_ram.sv:466:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:468:13
								initial begin
									// Trace: src/VX_dp_ram.sv:469:17
									begin : sv2v_autoblock_27
										// Trace: src/VX_dp_ram.sv:469:22
										integer i;
										// Trace: src/VX_dp_ram.sv:469:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:470:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:475:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:476:25
							if (write)
								// Trace: src/VX_dp_ram.sv:477:29
								ram[waddr] <= wdata;
						// Trace: src/VX_dp_ram.sv:480:21
						assign rdata = ram[raddr];
					end
				end
				else begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:484:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:487:13
								initial begin
									// Trace: src/VX_dp_ram.sv:487:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:489:13
								initial begin
									// Trace: src/VX_dp_ram.sv:490:17
									begin : sv2v_autoblock_28
										// Trace: src/VX_dp_ram.sv:490:22
										integer i;
										// Trace: src/VX_dp_ram.sv:490:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:491:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:496:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:497:25
							if (write)
								// Trace: src/VX_dp_ram.sv:498:29
								begin : sv2v_autoblock_29
									// Trace: src/VX_dp_ram.sv:498:34
									integer i;
									// Trace: src/VX_dp_ram.sv:498:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:499:33
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:500:37
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_dp_ram.sv:505:21
						assign rdata = ram[raddr];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:507:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:510:13
								initial begin
									// Trace: src/VX_dp_ram.sv:510:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:512:13
								initial begin
									// Trace: src/VX_dp_ram.sv:513:17
									begin : sv2v_autoblock_30
										// Trace: src/VX_dp_ram.sv:513:22
										integer i;
										// Trace: src/VX_dp_ram.sv:513:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:514:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:519:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:520:25
							if (write)
								// Trace: src/VX_dp_ram.sv:521:29
								ram[waddr] <= wdata;
						// Trace: src/VX_dp_ram.sv:524:21
						assign rdata = ram[raddr];
					end
				end
			end
		end
	endgenerate
endmodule
// removed module with interface ports: VX_csr_unit
module VX_cache_data (
	clk,
	reset,
	stall,
	init,
	fill,
	flush,
	read,
	write,
	line_idx,
	evict_way,
	tag_matches,
	fill_data,
	write_word,
	write_byteen,
	word_idx,
	way_idx_r,
	read_data,
	evict_byteen
);
	// Trace: src/VX_cache_data.sv:2:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_cache_data.sv:3:15
	parameter LINE_SIZE = 16;
	// Trace: src/VX_cache_data.sv:4:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_data.sv:5:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_data.sv:6:15
	parameter WORD_SIZE = 1;
	// Trace: src/VX_cache_data.sv:7:15
	parameter WRITE_ENABLE = 1;
	// Trace: src/VX_cache_data.sv:8:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_cache_data.sv:9:15
	parameter DIRTY_BYTES = 0;
	// Trace: src/VX_cache_data.sv:11:5
	input wire clk;
	// Trace: src/VX_cache_data.sv:12:5
	input wire reset;
	// Trace: src/VX_cache_data.sv:13:5
	input wire stall;
	// Trace: src/VX_cache_data.sv:14:5
	input wire init;
	// Trace: src/VX_cache_data.sv:15:5
	input wire fill;
	// Trace: src/VX_cache_data.sv:16:5
	input wire flush;
	// Trace: src/VX_cache_data.sv:17:5
	input wire read;
	// Trace: src/VX_cache_data.sv:18:5
	input wire write;
	// Trace: src/VX_cache_data.sv:19:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx;
	// Trace: src/VX_cache_data.sv:20:5
	input wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] evict_way;
	// Trace: src/VX_cache_data.sv:21:5
	input wire [NUM_WAYS - 1:0] tag_matches;
	// Trace: src/VX_cache_data.sv:22:5
	input wire [((LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] fill_data;
	// Trace: src/VX_cache_data.sv:23:5
	input wire [(8 * WORD_SIZE) - 1:0] write_word;
	// Trace: src/VX_cache_data.sv:24:5
	input wire [WORD_SIZE - 1:0] write_byteen;
	// Trace: src/VX_cache_data.sv:25:5
	input wire [($clog2(LINE_SIZE / WORD_SIZE) > 0 ? $clog2(LINE_SIZE / WORD_SIZE) : 1) - 1:0] word_idx;
	// Trace: src/VX_cache_data.sv:26:5
	input wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] way_idx_r;
	// Trace: src/VX_cache_data.sv:27:5
	output wire [(8 * LINE_SIZE) - 1:0] read_data;
	// Trace: src/VX_cache_data.sv:28:5
	output wire [LINE_SIZE - 1:0] evict_byteen;
	// Trace: src/VX_cache_data.sv:30:5
	wire [((LINE_SIZE / WORD_SIZE) * WORD_SIZE) - 1:0] write_mask;
	// Trace: src/VX_cache_data.sv:31:5
	genvar _gv_i_194;
	generate
		for (_gv_i_194 = 0; _gv_i_194 < (LINE_SIZE / WORD_SIZE); _gv_i_194 = _gv_i_194 + 1) begin : g_write_mask
			localparam i = _gv_i_194;
			// Trace: src/VX_cache_data.sv:32:9
			wire word_en = ((LINE_SIZE / WORD_SIZE) == 1) || (word_idx == i);
			// Trace: src/VX_cache_data.sv:33:9
			assign write_mask[i * WORD_SIZE+:WORD_SIZE] = write_byteen & {WORD_SIZE {word_en}};
		end
	endgenerate
	// Trace: src/VX_cache_data.sv:35:5
	generate
		if (DIRTY_BYTES != 0) begin : g_dirty_bytes
			// Trace: src/VX_cache_data.sv:36:9
			wire [(NUM_WAYS * LINE_SIZE) - 1:0] byteen_rdata;
			genvar _gv_i_195;
			for (_gv_i_195 = 0; _gv_i_195 < NUM_WAYS; _gv_i_195 = _gv_i_195 + 1) begin : g_byteen_store
				localparam i = _gv_i_195;
				// Trace: src/VX_cache_data.sv:38:13
				wire [LINE_SIZE - 1:0] byteen_wdata = {LINE_SIZE {write}};
				// Trace: src/VX_cache_data.sv:39:13
				wire [LINE_SIZE - 1:0] byteen_wren = {LINE_SIZE {(init || fill) || flush}} | write_mask;
				// Trace: src/VX_cache_data.sv:40:13
				wire byteen_write = (((fill || flush) && ((NUM_WAYS == 1) || (evict_way == i))) || (write && tag_matches[i])) || init;
				// Trace: src/VX_cache_data.sv:43:13
				wire byteen_read = fill || flush;
				// Trace: src/VX_cache_data.sv:44:13
				VX_sp_ram #(
					.DATAW(LINE_SIZE),
					.WRENW(LINE_SIZE),
					.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
					.OUT_REG(1),
					.RDW_MODE("R")
				) byteen_store(
					.clk(clk),
					.reset(reset),
					.read(byteen_read),
					.write(byteen_write),
					.wren(byteen_wren),
					.addr(line_idx),
					.wdata(byteen_wdata),
					.rdata(byteen_rdata[i * LINE_SIZE+:LINE_SIZE])
				);
			end
			// Trace: src/VX_cache_data.sv:61:9
			assign evict_byteen = byteen_rdata[way_idx_r * LINE_SIZE+:LINE_SIZE];
		end
		else begin : g_no_dirty_bytes
			// Trace: src/VX_cache_data.sv:63:9
			assign evict_byteen = 1'sb1;
		end
	endgenerate
	// Trace: src/VX_cache_data.sv:65:5
	wire [((NUM_WAYS * (LINE_SIZE / WORD_SIZE)) * (8 * WORD_SIZE)) - 1:0] line_rdata;
	// Trace: src/VX_cache_data.sv:66:5
	genvar _gv_i_196;
	generate
		for (_gv_i_196 = 0; _gv_i_196 < NUM_WAYS; _gv_i_196 = _gv_i_196 + 1) begin : g_data_store
			localparam i = _gv_i_196;
			// Trace: src/VX_cache_data.sv:67:9
			localparam WRENW = (WRITE_ENABLE ? LINE_SIZE : 1);
			// Trace: src/VX_cache_data.sv:68:9
			wire [((LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] line_wdata;
			// Trace: src/VX_cache_data.sv:69:9
			wire [WRENW - 1:0] line_wren;
			if (WRITE_ENABLE) begin : g_wren
				// Trace: src/VX_cache_data.sv:71:13
				assign line_wdata = (fill ? fill_data : {LINE_SIZE / WORD_SIZE {write_word}});
				// Trace: src/VX_cache_data.sv:72:13
				assign line_wren = {LINE_SIZE {fill}} | write_mask;
			end
			else begin : g_no_wren
				// Trace: src/VX_cache_data.sv:74:13
				assign line_wdata = fill_data;
				// Trace: src/VX_cache_data.sv:75:13
				assign line_wren = 1'b1;
			end
			// Trace: src/VX_cache_data.sv:77:9
			wire line_write = (fill && ((NUM_WAYS == 1) || (evict_way == i))) || ((write && tag_matches[i]) && WRITE_ENABLE);
			// Trace: src/VX_cache_data.sv:79:9
			wire line_read = read || ((fill || flush) && WRITEBACK);
			// Trace: src/VX_cache_data.sv:80:9
			VX_sp_ram #(
				.DATAW(8 * LINE_SIZE),
				.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
				.WRENW(WRENW),
				.OUT_REG(1),
				.RDW_MODE("R")
			) data_store(
				.clk(clk),
				.reset(reset),
				.read(line_read),
				.write(line_write),
				.wren(line_wren),
				.addr(line_idx),
				.wdata(line_wdata),
				.rdata(line_rdata[(8 * WORD_SIZE) * (i * (LINE_SIZE / WORD_SIZE))+:(8 * WORD_SIZE) * (LINE_SIZE / WORD_SIZE)])
			);
		end
	endgenerate
	// Trace: src/VX_cache_data.sv:97:5
	assign read_data = line_rdata[(8 * WORD_SIZE) * (way_idx_r * (LINE_SIZE / WORD_SIZE))+:(8 * WORD_SIZE) * (LINE_SIZE / WORD_SIZE)];
endmodule
module VX_rr_arbiter (
	clk,
	reset,
	requests,
	grant_index,
	grant_onehot,
	grant_valid,
	grant_ready
);
	// Trace: src/VX_rr_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_rr_arbiter.sv:3:15
	parameter MODEL = 1;
	// Trace: src/VX_rr_arbiter.sv:4:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_rr_arbiter.sv:5:15
	parameter LUT_OPT = 0;
	// Trace: src/VX_rr_arbiter.sv:7:5
	input wire clk;
	// Trace: src/VX_rr_arbiter.sv:8:5
	input wire reset;
	// Trace: src/VX_rr_arbiter.sv:9:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_rr_arbiter.sv:10:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_rr_arbiter.sv:11:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_rr_arbiter.sv:12:5
	output wire grant_valid;
	// Trace: src/VX_rr_arbiter.sv:13:5
	input wire grant_ready;
	// Trace: src/VX_rr_arbiter.sv:15:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_REQS == 1) begin : g_passthru
			// Trace: src/VX_rr_arbiter.sv:16:9
			assign grant_index = 1'sb0;
			// Trace: src/VX_rr_arbiter.sv:17:9
			assign grant_onehot = requests;
			// Trace: src/VX_rr_arbiter.sv:18:9
			assign grant_valid = requests[0];
		end
		else if (LUT_OPT && (NUM_REQS == 2)) begin : g_lut2
			// Trace: src/VX_rr_arbiter.sv:20:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:21:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:22:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:23:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:24:13
				casez ({state, requests})
					3'b001, 3'b1z1: begin
						// Trace: src/VX_rr_arbiter.sv:26:28
						grant_onehot_w = 2'b01;
						// Trace: src/VX_rr_arbiter.sv:26:52
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					3'b01z, 3'b110: begin
						// Trace: src/VX_rr_arbiter.sv:28:28
						grant_onehot_w = 2'b10;
						// Trace: src/VX_rr_arbiter.sv:28:52
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:29:28
						grant_onehot_w = 2'b00;
						// Trace: src/VX_rr_arbiter.sv:29:52
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:32:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:33:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:34:17
					state <= 1'sb0;
				else if (grant_ready)
					// Trace: src/VX_rr_arbiter.sv:36:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:39:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:40:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:41:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 3)) begin : g_lut3
			// Trace: src/VX_rr_arbiter.sv:43:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:44:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:45:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:46:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:47:13
				casez ({state, requests})
					5'b00001, 5'b010z1, 5'b10zz1: begin
						// Trace: src/VX_rr_arbiter.sv:50:30
						grant_onehot_w = 3'b001;
						// Trace: src/VX_rr_arbiter.sv:50:55
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					5'b00z1z, 5'b01010, 5'b10z10: begin
						// Trace: src/VX_rr_arbiter.sv:53:30
						grant_onehot_w = 3'b010;
						// Trace: src/VX_rr_arbiter.sv:53:55
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					5'b0010z, 5'b011zz, 5'b10100: begin
						// Trace: src/VX_rr_arbiter.sv:56:30
						grant_onehot_w = 3'b100;
						// Trace: src/VX_rr_arbiter.sv:56:55
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:57:30
						grant_onehot_w = 3'b000;
						// Trace: src/VX_rr_arbiter.sv:57:55
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:60:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:61:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:62:17
					state <= 1'sb0;
				else if (grant_ready)
					// Trace: src/VX_rr_arbiter.sv:64:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:67:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:68:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:69:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 4)) begin : g_lut4
			// Trace: src/VX_rr_arbiter.sv:71:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:72:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:73:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:74:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:75:13
				casez ({state, requests})
					6'b000001, 6'b0100z1, 6'b100zz1, 6'b11zzz1: begin
						// Trace: src/VX_rr_arbiter.sv:79:31
						grant_onehot_w = 4'b0001;
						// Trace: src/VX_rr_arbiter.sv:79:57
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					6'b00zz1z, 6'b010010, 6'b100z10, 6'b11zz10: begin
						// Trace: src/VX_rr_arbiter.sv:83:31
						grant_onehot_w = 4'b0010;
						// Trace: src/VX_rr_arbiter.sv:83:57
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					6'b00z10z, 6'b01z1zz, 6'b100100, 6'b11z100: begin
						// Trace: src/VX_rr_arbiter.sv:87:31
						grant_onehot_w = 4'b0100;
						// Trace: src/VX_rr_arbiter.sv:87:57
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					6'b00100z, 6'b0110zz, 6'b101zzz, 6'b111000: begin
						// Trace: src/VX_rr_arbiter.sv:91:31
						grant_onehot_w = 4'b1000;
						// Trace: src/VX_rr_arbiter.sv:91:57
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:92:31
						grant_onehot_w = 4'b0000;
						// Trace: src/VX_rr_arbiter.sv:92:57
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:95:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:96:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:97:17
					state <= 1'sb0;
				else if (grant_ready)
					// Trace: src/VX_rr_arbiter.sv:99:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:102:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:103:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:104:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 5)) begin : g_lut5
			// Trace: src/VX_rr_arbiter.sv:106:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:107:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:108:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:109:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:110:13
				casez ({state, requests})
					8'b00000001, 8'b001000z1, 8'b01000zz1, 8'b0110zzz1, 8'b100zzzz1: begin
						// Trace: src/VX_rr_arbiter.sv:115:33
						grant_onehot_w = 5'b00001;
						// Trace: src/VX_rr_arbiter.sv:115:60
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					8'b000zzz1z, 8'b00100010, 8'b01000z10, 8'b0110zz10, 8'b100zzz10: begin
						// Trace: src/VX_rr_arbiter.sv:120:33
						grant_onehot_w = 5'b00010;
						// Trace: src/VX_rr_arbiter.sv:120:60
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					8'b000zz10z, 8'b001zz1zz, 8'b01000100, 8'b0110z100, 8'b100zz100: begin
						// Trace: src/VX_rr_arbiter.sv:125:33
						grant_onehot_w = 5'b00100;
						// Trace: src/VX_rr_arbiter.sv:125:60
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					8'b000z100z, 8'b001z10zz, 8'b010z1zzz, 8'b01101000, 8'b100z1000: begin
						// Trace: src/VX_rr_arbiter.sv:130:33
						grant_onehot_w = 5'b01000;
						// Trace: src/VX_rr_arbiter.sv:130:60
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					8'b0001000z, 8'b001100zz, 8'b01010zzz, 8'b0111zzzz, 8'b10010000: begin
						// Trace: src/VX_rr_arbiter.sv:135:33
						grant_onehot_w = 5'b10000;
						// Trace: src/VX_rr_arbiter.sv:135:60
						grant_index_w = sv2v_cast_76B5F_signed(4);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:136:33
						grant_onehot_w = 5'b00000;
						// Trace: src/VX_rr_arbiter.sv:136:60
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:139:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:140:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:141:17
					state <= 1'sb0;
				else if (grant_ready)
					// Trace: src/VX_rr_arbiter.sv:143:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:146:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:147:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:148:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 6)) begin : g_lut6
			// Trace: src/VX_rr_arbiter.sv:150:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:151:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:152:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:153:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:154:13
				casez ({state, requests})
					9'b000000001, 9'b0010000z1, 9'b010000zz1, 9'b01100zzz1, 9'b1000zzzz1, 9'b101zzzzz1: begin
						// Trace: src/VX_rr_arbiter.sv:160:34
						grant_onehot_w = 6'b000001;
						// Trace: src/VX_rr_arbiter.sv:160:62
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					9'b000zzzz1z, 9'b001000010, 9'b010000z10, 9'b01100zz10, 9'b1000zzz10, 9'b101zzzz10: begin
						// Trace: src/VX_rr_arbiter.sv:166:34
						grant_onehot_w = 6'b000010;
						// Trace: src/VX_rr_arbiter.sv:166:62
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					9'b000zzz10z, 9'b001zzz1zz, 9'b010000100, 9'b01100z100, 9'b1000zz100, 9'b101zzz100: begin
						// Trace: src/VX_rr_arbiter.sv:172:34
						grant_onehot_w = 6'b000100;
						// Trace: src/VX_rr_arbiter.sv:172:62
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					9'b000zz100z, 9'b001zz10zz, 9'b010zz1zzz, 9'b011001000, 9'b1000z1000, 9'b101zz1000: begin
						// Trace: src/VX_rr_arbiter.sv:178:34
						grant_onehot_w = 6'b001000;
						// Trace: src/VX_rr_arbiter.sv:178:62
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					9'b000z1000z, 9'b001z100zz, 9'b010z10zzz, 9'b011z1zzzz, 9'b100010000, 9'b101z10000: begin
						// Trace: src/VX_rr_arbiter.sv:184:34
						grant_onehot_w = 6'b010000;
						// Trace: src/VX_rr_arbiter.sv:184:62
						grant_index_w = sv2v_cast_76B5F_signed(4);
					end
					9'b00010000z, 9'b0011000zz, 9'b010100zzz, 9'b01110zzzz, 9'b1001zzzzz, 9'b101100000: begin
						// Trace: src/VX_rr_arbiter.sv:190:34
						grant_onehot_w = 6'b100000;
						// Trace: src/VX_rr_arbiter.sv:190:62
						grant_index_w = sv2v_cast_76B5F_signed(5);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:191:34
						grant_onehot_w = 6'b000000;
						// Trace: src/VX_rr_arbiter.sv:191:62
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:194:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:195:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:196:17
					state <= 1'sb0;
				else if (grant_ready)
					// Trace: src/VX_rr_arbiter.sv:198:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:201:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:202:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:203:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 7)) begin : g_lut7
			// Trace: src/VX_rr_arbiter.sv:205:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:206:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:207:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:208:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:209:13
				casez ({state, requests})
					10'b0000000001, 10'b00100000z1, 10'b0100000zz1, 10'b011000zzz1, 10'b100000zzz1, 10'b10100zzzz1, 10'b110zzzzzz1: begin
						// Trace: src/VX_rr_arbiter.sv:216:36
						grant_onehot_w = 7'b0000001;
						// Trace: src/VX_rr_arbiter.sv:216:65
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					10'b000zzzzz1z, 10'b0010000010, 10'b0100000z10, 10'b011000zz10, 10'b10000zzz10, 10'b1010zzzz10, 10'b110zzzzz10: begin
						// Trace: src/VX_rr_arbiter.sv:223:36
						grant_onehot_w = 7'b0000010;
						// Trace: src/VX_rr_arbiter.sv:223:65
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					10'b000zzzz10z, 10'b001zzzz1zz, 10'b0100000100, 10'b011000z100, 10'b10000zz100, 10'b1010zzz100, 10'b110zzzz100: begin
						// Trace: src/VX_rr_arbiter.sv:230:36
						grant_onehot_w = 7'b0000100;
						// Trace: src/VX_rr_arbiter.sv:230:65
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					10'b000zzz100z, 10'b001zzz10zz, 10'b010zzz1zzz, 10'b0110001000, 10'b10000z1000, 10'b1010zz1000, 10'b110zzz1000: begin
						// Trace: src/VX_rr_arbiter.sv:237:36
						grant_onehot_w = 7'b0001000;
						// Trace: src/VX_rr_arbiter.sv:237:65
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					10'b000zz1000z, 10'b001zz100zz, 10'b010zz10zzz, 10'b011zz1zzzz, 10'b1000010000, 10'b1010z10000, 10'b110zz10000: begin
						// Trace: src/VX_rr_arbiter.sv:244:36
						grant_onehot_w = 7'b0010000;
						// Trace: src/VX_rr_arbiter.sv:244:65
						grant_index_w = sv2v_cast_76B5F_signed(4);
					end
					10'b000z10000z, 10'b001z1000zz, 10'b010z100zzz, 10'b011z10zzzz, 10'b100z1zzzzz, 10'b1010100000, 10'b110z100000: begin
						// Trace: src/VX_rr_arbiter.sv:251:36
						grant_onehot_w = 7'b0100000;
						// Trace: src/VX_rr_arbiter.sv:251:65
						grant_index_w = sv2v_cast_76B5F_signed(5);
					end
					10'b000100000z, 10'b00110000zz, 10'b0101000zzz, 10'b011100zzzz, 10'b10010zzzzz, 10'b1011zzzzzz, 10'b1101000000: begin
						// Trace: src/VX_rr_arbiter.sv:258:36
						grant_onehot_w = 7'b1000000;
						// Trace: src/VX_rr_arbiter.sv:258:65
						grant_index_w = sv2v_cast_76B5F_signed(6);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:259:35
						grant_onehot_w = 7'b0000000;
						// Trace: src/VX_rr_arbiter.sv:259:64
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:262:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:263:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:264:17
					state <= 1'sb0;
				else if (grant_ready)
					// Trace: src/VX_rr_arbiter.sv:266:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:269:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:270:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:271:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 8)) begin : g_lut8
			// Trace: src/VX_rr_arbiter.sv:273:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:274:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:275:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:276:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:277:13
				casez ({state, requests})
					11'b00000000001, 11'b001000000z1, 11'b01000000zz1, 11'b0110000zzz1, 11'b100000zzzz1, 11'b10100zzzzz1, 11'b1100zzzzzz1, 11'b111zzzzzzz1: begin
						// Trace: src/VX_rr_arbiter.sv:285:37
						grant_onehot_w = 8'b00000001;
						// Trace: src/VX_rr_arbiter.sv:285:67
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					11'b000zzzzzz1z, 11'b00100000010, 11'b01000000z10, 11'b0110000zz10, 11'b100000zzz10, 11'b10100zzzz10, 11'b1100zzzzz10, 11'b111zzzzzz10: begin
						// Trace: src/VX_rr_arbiter.sv:293:37
						grant_onehot_w = 8'b00000010;
						// Trace: src/VX_rr_arbiter.sv:293:67
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					11'b000zzzzz10z, 11'b001zzzzz1zz, 11'b01000000100, 11'b0110000z100, 11'b100000zz100, 11'b10100zzz100, 11'b1100zzzz100, 11'b111zzzzz100: begin
						// Trace: src/VX_rr_arbiter.sv:301:37
						grant_onehot_w = 8'b00000100;
						// Trace: src/VX_rr_arbiter.sv:301:67
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					11'b000zzzz100z, 11'b001zzzz10zz, 11'b010zzzz1zzz, 11'b01100001000, 11'b100000z1000, 11'b10100zz1000, 11'b1100zzz1000, 11'b111zzzz1000: begin
						// Trace: src/VX_rr_arbiter.sv:309:37
						grant_onehot_w = 8'b00001000;
						// Trace: src/VX_rr_arbiter.sv:309:67
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					11'b000zzz1000z, 11'b001zzz100zz, 11'b010zzz10zzz, 11'b011zzz1zzzz, 11'b10000010000, 11'b10100z10000, 11'b1100zz10000, 11'b111zzz10000: begin
						// Trace: src/VX_rr_arbiter.sv:317:37
						grant_onehot_w = 8'b00010000;
						// Trace: src/VX_rr_arbiter.sv:317:67
						grant_index_w = sv2v_cast_76B5F_signed(4);
					end
					11'b000zz10000z, 11'b001zz1000zz, 11'b010zz100zzz, 11'b011zz10zzzz, 11'b100zz1zzzzz, 11'b10100100000, 11'b1100z100000, 11'b111zz100000: begin
						// Trace: src/VX_rr_arbiter.sv:325:37
						grant_onehot_w = 8'b00100000;
						// Trace: src/VX_rr_arbiter.sv:325:67
						grant_index_w = sv2v_cast_76B5F_signed(5);
					end
					11'b000z100000z, 11'b001z10000zz, 11'b010z1000zzz, 11'b011z100zzzz, 11'b100z10zzzzz, 11'b101z1zzzzzz, 11'b11001000000, 11'b111z1000000: begin
						// Trace: src/VX_rr_arbiter.sv:333:37
						grant_onehot_w = 8'b01000000;
						// Trace: src/VX_rr_arbiter.sv:333:67
						grant_index_w = sv2v_cast_76B5F_signed(6);
					end
					11'b0001000000z, 11'b001100000zz, 11'b01010000zzz, 11'b0111000zzzz, 11'b100100zzzzz, 11'b10110zzzzzz, 11'b1101zzzzzzz, 11'b11110000000: begin
						// Trace: src/VX_rr_arbiter.sv:341:37
						grant_onehot_w = 8'b10000000;
						// Trace: src/VX_rr_arbiter.sv:341:67
						grant_index_w = sv2v_cast_76B5F_signed(7);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:342:37
						grant_onehot_w = 8'b00000000;
						// Trace: src/VX_rr_arbiter.sv:342:67
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:345:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:346:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:347:17
					state <= 1'sb0;
				else if (grant_ready)
					// Trace: src/VX_rr_arbiter.sv:349:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:352:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:353:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:354:9
			assign grant_valid = |requests;
		end
		else if (MODEL == 1) begin : g_model1
			// Trace: src/VX_rr_arbiter.sv:356:9
			wire [NUM_REQS - 1:0] masked_pri_reqs;
			wire [NUM_REQS - 1:0] unmasked_pri_reqs;
			// Trace: src/VX_rr_arbiter.sv:357:9
			reg [NUM_REQS - 1:0] reqs_mask;
			// Trace: src/VX_rr_arbiter.sv:358:9
			wire [NUM_REQS - 1:0] masked_reqs = requests & reqs_mask;
			// Trace: src/VX_rr_arbiter.sv:359:9
			assign masked_pri_reqs[0] = 1'b0;
			genvar _gv_i_197;
			for (_gv_i_197 = 1; _gv_i_197 < NUM_REQS; _gv_i_197 = _gv_i_197 + 1) begin : g_masked_pri_reqs
				localparam i = _gv_i_197;
				// Trace: src/VX_rr_arbiter.sv:361:13
				assign masked_pri_reqs[i] = masked_pri_reqs[i - 1] | masked_reqs[i - 1];
			end
			// Trace: src/VX_rr_arbiter.sv:363:9
			assign unmasked_pri_reqs[0] = 1'b0;
			genvar _gv_i_198;
			for (_gv_i_198 = 1; _gv_i_198 < NUM_REQS; _gv_i_198 = _gv_i_198 + 1) begin : g_unmasked_pri_reqs
				localparam i = _gv_i_198;
				// Trace: src/VX_rr_arbiter.sv:365:13
				assign unmasked_pri_reqs[i] = unmasked_pri_reqs[i - 1] | requests[i - 1];
			end
			// Trace: src/VX_rr_arbiter.sv:367:9
			wire [NUM_REQS - 1:0] grant_masked = masked_reqs & ~masked_pri_reqs;
			// Trace: src/VX_rr_arbiter.sv:368:9
			wire [NUM_REQS - 1:0] grant_unmasked = requests & ~unmasked_pri_reqs;
			// Trace: src/VX_rr_arbiter.sv:369:9
			wire has_masked_reqs = |masked_reqs;
			// Trace: src/VX_rr_arbiter.sv:370:9
			wire has_unmasked_reqs = |requests;
			// Trace: src/VX_rr_arbiter.sv:371:9
			assign grant_onehot = (has_masked_reqs ? grant_masked : grant_unmasked);
			// Trace: src/VX_rr_arbiter.sv:372:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:373:7
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:374:5
					reqs_mask <= {NUM_REQS {1'b1}};
				else if (grant_ready) begin
					begin
						// Trace: src/VX_rr_arbiter.sv:376:5
						if (has_masked_reqs)
							// Trace: src/VX_rr_arbiter.sv:377:21
							reqs_mask <= masked_pri_reqs;
						else if (has_unmasked_reqs)
							// Trace: src/VX_rr_arbiter.sv:379:21
							reqs_mask <= unmasked_pri_reqs;
					end
				end
			// Trace: src/VX_rr_arbiter.sv:383:9
			VX_onehot_encoder #(.N(NUM_REQS)) onehot_encoder(
				.data_in(grant_onehot),
				.data_out(grant_index),
				.valid_out(grant_valid)
			);
		end
		else if (MODEL == 2) begin : g_model2
			// Trace: src/VX_rr_arbiter.sv:391:9
			reg [(NUM_REQS * LOG_NUM_REQS) - 1:0] grant_table;
			// Trace: src/VX_rr_arbiter.sv:392:9
			reg [LOG_NUM_REQS - 1:0] state;
			genvar _gv_i_199;
			for (_gv_i_199 = 0; _gv_i_199 < NUM_REQS; _gv_i_199 = _gv_i_199 + 1) begin : g_grant_table
				localparam i = _gv_i_199;
				// Trace: src/VX_rr_arbiter.sv:394:13
				always @(*) begin
					// Trace: src/VX_rr_arbiter.sv:395:17
					grant_table[i * LOG_NUM_REQS+:LOG_NUM_REQS] = 1'sbx;
					// Trace: src/VX_rr_arbiter.sv:396:17
					begin : sv2v_autoblock_1
						// Trace: src/VX_rr_arbiter.sv:396:22
						integer j;
						// Trace: src/VX_rr_arbiter.sv:396:22
						for (j = NUM_REQS - 1; j >= 0; j = j - 1)
							begin
								// Trace: src/VX_rr_arbiter.sv:397:21
								if (requests[((i + j) + 1) % NUM_REQS])
									// Trace: src/VX_rr_arbiter.sv:398:25
									grant_table[i * LOG_NUM_REQS+:LOG_NUM_REQS] = sv2v_cast_76B5F_signed(((i + j) + 1) % NUM_REQS);
							end
					end
				end
			end
			// Trace: src/VX_rr_arbiter.sv:403:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:404:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:405:17
					state <= 0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:407:17
					state <= grant_index;
			// Trace: src/VX_rr_arbiter.sv:410:9
			VX_demux #(
				.DATAW(1),
				.N(NUM_REQS)
			) grant_decoder(
				.sel_in(grant_index),
				.data_in(grant_valid),
				.data_out(grant_onehot)
			);
			// Trace: src/VX_rr_arbiter.sv:418:9
			assign grant_index = grant_table[state * LOG_NUM_REQS+:LOG_NUM_REQS];
			// Trace: src/VX_rr_arbiter.sv:419:9
			assign grant_valid = |requests;
		end
	endgenerate
endmodule
// removed interface: VX_writeback_if
// removed module with interface ports: VX_alu_unit
// removed module with interface ports: VX_mem_unit
// removed interface: VX_commit_if
// removed module with interface ports: VX_gather_unit
// removed module with interface ports: VX_cluster
module VX_find_first (
	data_in,
	valid_in,
	data_out,
	valid_out
);
	// Trace: src/VX_find_first.sv:2:15
	parameter N = 1;
	// Trace: src/VX_find_first.sv:3:15
	parameter DATAW = 1;
	// Trace: src/VX_find_first.sv:4:15
	parameter REVERSE = 0;
	// Trace: src/VX_find_first.sv:6:5
	input wire [(N * DATAW) - 1:0] data_in;
	// Trace: src/VX_find_first.sv:7:5
	input wire [N - 1:0] valid_in;
	// Trace: src/VX_find_first.sv:8:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_find_first.sv:9:5
	output wire valid_out;
	// Trace: src/VX_find_first.sv:11:5
	localparam LOGN = $clog2(N);
	// Trace: src/VX_find_first.sv:12:5
	localparam TL = (1 << LOGN) - 1;
	// Trace: src/VX_find_first.sv:13:5
	localparam TN = (1 << (LOGN + 1)) - 1;
	// Trace: src/VX_find_first.sv:14:5
	wire s_n [0:TN - 1];
	// Trace: src/VX_find_first.sv:15:5
	wire [DATAW - 1:0] d_n [0:TN - 1];
	// Trace: src/VX_find_first.sv:16:5
	genvar _gv_i_211;
	generate
		for (_gv_i_211 = 0; _gv_i_211 < N; _gv_i_211 = _gv_i_211 + 1) begin : g_reverse
			localparam i = _gv_i_211;
			// Trace: src/VX_find_first.sv:17:9
			assign s_n[TL + i] = (REVERSE ? valid_in[(N - 1) - i] : valid_in[i]);
			// Trace: src/VX_find_first.sv:18:9
			assign d_n[TL + i] = (REVERSE ? data_in[((N - 1) - i) * DATAW+:DATAW] : data_in[i * DATAW+:DATAW]);
		end
	endgenerate
	// Trace: src/VX_find_first.sv:20:5
	generate
		if (TL < (TN - N)) begin : g_fill
			genvar _gv_i_212;
			for (_gv_i_212 = TL + N; _gv_i_212 < TN; _gv_i_212 = _gv_i_212 + 1) begin : g_i
				localparam i = _gv_i_212;
				// Trace: src/VX_find_first.sv:22:13
				assign s_n[i] = 0;
				// Trace: src/VX_find_first.sv:23:13
				assign d_n[i] = 1'sb0;
			end
		end
	endgenerate
	// Trace: src/VX_find_first.sv:26:5
	genvar _gv_j_22;
	generate
		for (_gv_j_22 = 0; _gv_j_22 < LOGN; _gv_j_22 = _gv_j_22 + 1) begin : g_scan
			localparam j = _gv_j_22;
			// Trace: src/VX_find_first.sv:27:9
			localparam I = 1 << j;
			genvar _gv_i_213;
			for (_gv_i_213 = 0; _gv_i_213 < I; _gv_i_213 = _gv_i_213 + 1) begin : g_i
				localparam i = _gv_i_213;
				// Trace: src/VX_find_first.sv:29:13
				localparam K = (I + i) - 1;
				// Trace: src/VX_find_first.sv:30:13
				assign s_n[K] = s_n[(2 * K) + 1] | s_n[(2 * K) + 2];
				// Trace: src/VX_find_first.sv:31:13
				assign d_n[K] = (s_n[(2 * K) + 1] ? d_n[(2 * K) + 1] : d_n[(2 * K) + 2]);
			end
		end
	endgenerate
	// Trace: src/VX_find_first.sv:34:5
	assign valid_out = s_n[0];
	// Trace: src/VX_find_first.sv:35:5
	assign data_out = d_n[0];
endmodule
module VX_sp_ram (
	clk,
	reset,
	read,
	write,
	wren,
	addr,
	wdata,
	rdata
);
	// Trace: src/VX_sp_ram.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_sp_ram.sv:3:15
	parameter SIZE = 1;
	// Trace: src/VX_sp_ram.sv:4:15
	parameter WRENW = 1;
	// Trace: src/VX_sp_ram.sv:5:15
	parameter OUT_REG = 0;
	// Trace: src/VX_sp_ram.sv:6:15
	parameter LUTRAM = 0;
	// Trace: src/VX_sp_ram.sv:7:15
	parameter RDW_MODE = "W";
	// Trace: src/VX_sp_ram.sv:8:15
	parameter RADDR_REG = 0;
	// Trace: src/VX_sp_ram.sv:9:15
	parameter RDW_ASSERT = 0;
	// Trace: src/VX_sp_ram.sv:10:15
	parameter RESET_RAM = 0;
	// Trace: src/VX_sp_ram.sv:11:15
	parameter INIT_ENABLE = 0;
	// Trace: src/VX_sp_ram.sv:12:15
	parameter INIT_FILE = "";
	// Trace: src/VX_sp_ram.sv:13:15
	parameter [DATAW - 1:0] INIT_VALUE = 0;
	// Trace: src/VX_sp_ram.sv:14:15
	parameter ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
	// Trace: src/VX_sp_ram.sv:16:5
	input wire clk;
	// Trace: src/VX_sp_ram.sv:17:5
	input wire reset;
	// Trace: src/VX_sp_ram.sv:18:5
	input wire read;
	// Trace: src/VX_sp_ram.sv:19:5
	input wire write;
	// Trace: src/VX_sp_ram.sv:20:5
	input wire [WRENW - 1:0] wren;
	// Trace: src/VX_sp_ram.sv:21:5
	input wire [ADDRW - 1:0] addr;
	// Trace: src/VX_sp_ram.sv:22:5
	input wire [DATAW - 1:0] wdata;
	// Trace: src/VX_sp_ram.sv:23:5
	output wire [DATAW - 1:0] rdata;
	// Trace: src/VX_sp_ram.sv:25:5
	localparam WSELW = DATAW / WRENW;
	// Trace: src/VX_sp_ram.sv:26:5
	localparam FORCE_BRAM = !LUTRAM && ((SIZE * DATAW) >= 1024);
	// Trace: src/VX_sp_ram.sv:27:5
	generate
		if (OUT_REG) begin : g_sync
			if (FORCE_BRAM) begin : g_bram
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:31:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:34:13
								initial begin
									// Trace: src/VX_sp_ram.sv:34:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:36:13
								initial begin
									// Trace: src/VX_sp_ram.sv:37:17
									begin : sv2v_autoblock_1
										// Trace: src/VX_sp_ram.sv:37:22
										integer i;
										// Trace: src/VX_sp_ram.sv:37:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:38:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:43:21
						reg [ADDRW - 1:0] addr_r;
						// Trace: src/VX_sp_ram.sv:44:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:45:25
							if (read || write) begin
								// Trace: src/VX_sp_ram.sv:46:29
								if (write)
									// Trace: src/VX_sp_ram.sv:47:33
									begin : sv2v_autoblock_2
										// Trace: src/VX_sp_ram.sv:47:38
										integer i;
										// Trace: src/VX_sp_ram.sv:47:38
										for (i = 0; i < WRENW; i = i + 1)
											begin
												// Trace: src/VX_sp_ram.sv:48:33
												if (wren[i])
													// Trace: src/VX_sp_ram.sv:49:37
													ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
											end
									end
								// Trace: src/VX_sp_ram.sv:53:29
								addr_r <= addr;
							end
						// Trace: src/VX_sp_ram.sv:56:21
						assign rdata = ram[addr_r];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:58:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:61:13
								initial begin
									// Trace: src/VX_sp_ram.sv:61:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:63:13
								initial begin
									// Trace: src/VX_sp_ram.sv:64:17
									begin : sv2v_autoblock_3
										// Trace: src/VX_sp_ram.sv:64:22
										integer i;
										// Trace: src/VX_sp_ram.sv:64:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:65:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:70:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:71:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:72:25
							if (read || write) begin
								begin
									// Trace: src/VX_sp_ram.sv:73:29
									if (write) begin
										// Trace: src/VX_sp_ram.sv:74:33
										ram[addr] <= wdata;
										// Trace: src/VX_sp_ram.sv:75:33
										rdata_r <= wdata;
									end
									else
										// Trace: src/VX_sp_ram.sv:77:33
										rdata_r <= ram[addr];
								end
							end
						// Trace: src/VX_sp_ram.sv:81:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "R") begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:85:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:88:13
								initial begin
									// Trace: src/VX_sp_ram.sv:88:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:90:13
								initial begin
									// Trace: src/VX_sp_ram.sv:91:17
									begin : sv2v_autoblock_4
										// Trace: src/VX_sp_ram.sv:91:22
										integer i;
										// Trace: src/VX_sp_ram.sv:91:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:92:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:97:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:98:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:99:25
							if (read || write) begin
								// Trace: src/VX_sp_ram.sv:100:29
								if (write)
									// Trace: src/VX_sp_ram.sv:101:33
									begin : sv2v_autoblock_5
										// Trace: src/VX_sp_ram.sv:101:38
										integer i;
										// Trace: src/VX_sp_ram.sv:101:38
										for (i = 0; i < WRENW; i = i + 1)
											begin
												// Trace: src/VX_sp_ram.sv:102:33
												if (wren[i])
													// Trace: src/VX_sp_ram.sv:103:37
													ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
											end
									end
								// Trace: src/VX_sp_ram.sv:107:29
								rdata_r <= ram[addr];
							end
						// Trace: src/VX_sp_ram.sv:110:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:112:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:115:13
								initial begin
									// Trace: src/VX_sp_ram.sv:115:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:117:13
								initial begin
									// Trace: src/VX_sp_ram.sv:118:17
									begin : sv2v_autoblock_6
										// Trace: src/VX_sp_ram.sv:118:22
										integer i;
										// Trace: src/VX_sp_ram.sv:118:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:119:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:124:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:125:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:126:25
							if (read || write) begin
								// Trace: src/VX_sp_ram.sv:127:29
								if (write)
									// Trace: src/VX_sp_ram.sv:128:33
									ram[addr] <= wdata;
								// Trace: src/VX_sp_ram.sv:130:29
								rdata_r <= ram[addr];
							end
						// Trace: src/VX_sp_ram.sv:133:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "N") begin : g_no_change
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:137:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:140:13
								initial begin
									// Trace: src/VX_sp_ram.sv:140:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:142:13
								initial begin
									// Trace: src/VX_sp_ram.sv:143:17
									begin : sv2v_autoblock_7
										// Trace: src/VX_sp_ram.sv:143:22
										integer i;
										// Trace: src/VX_sp_ram.sv:143:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:144:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:149:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:150:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:151:25
							if (read || write) begin
								begin
									// Trace: src/VX_sp_ram.sv:152:29
									if (write)
										// Trace: src/VX_sp_ram.sv:153:33
										begin : sv2v_autoblock_8
											// Trace: src/VX_sp_ram.sv:153:38
											integer i;
											// Trace: src/VX_sp_ram.sv:153:38
											for (i = 0; i < WRENW; i = i + 1)
												begin
													// Trace: src/VX_sp_ram.sv:154:33
													if (wren[i])
														// Trace: src/VX_sp_ram.sv:155:37
														ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
												end
										end
									else
										// Trace: src/VX_sp_ram.sv:159:33
										rdata_r <= ram[addr];
								end
							end
						// Trace: src/VX_sp_ram.sv:163:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:165:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:168:13
								initial begin
									// Trace: src/VX_sp_ram.sv:168:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:170:13
								initial begin
									// Trace: src/VX_sp_ram.sv:171:17
									begin : sv2v_autoblock_9
										// Trace: src/VX_sp_ram.sv:171:22
										integer i;
										// Trace: src/VX_sp_ram.sv:171:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:172:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:177:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:178:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:179:25
							if (read || write) begin
								begin
									// Trace: src/VX_sp_ram.sv:180:29
									if (write)
										// Trace: src/VX_sp_ram.sv:181:33
										ram[addr] <= wdata;
									else
										// Trace: src/VX_sp_ram.sv:183:33
										rdata_r <= ram[addr];
								end
							end
						// Trace: src/VX_sp_ram.sv:187:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "U") begin : g_undefined
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:191:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:194:13
								initial begin
									// Trace: src/VX_sp_ram.sv:194:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:196:13
								initial begin
									// Trace: src/VX_sp_ram.sv:197:17
									begin : sv2v_autoblock_10
										// Trace: src/VX_sp_ram.sv:197:22
										integer i;
										// Trace: src/VX_sp_ram.sv:197:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:198:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:203:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:204:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:205:25
							if (write)
								// Trace: src/VX_sp_ram.sv:206:29
								begin : sv2v_autoblock_11
									// Trace: src/VX_sp_ram.sv:206:34
									integer i;
									// Trace: src/VX_sp_ram.sv:206:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:207:33
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:208:37
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_sp_ram.sv:213:29
								rdata_r <= ram[addr];
						end
						// Trace: src/VX_sp_ram.sv:216:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:218:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:221:13
								initial begin
									// Trace: src/VX_sp_ram.sv:221:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:223:13
								initial begin
									// Trace: src/VX_sp_ram.sv:224:17
									begin : sv2v_autoblock_12
										// Trace: src/VX_sp_ram.sv:224:22
										integer i;
										// Trace: src/VX_sp_ram.sv:224:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:225:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:230:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:231:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:232:25
							if (write)
								// Trace: src/VX_sp_ram.sv:233:29
								ram[addr] <= wdata;
							if (read)
								// Trace: src/VX_sp_ram.sv:236:29
								rdata_r <= ram[addr];
						end
						// Trace: src/VX_sp_ram.sv:239:21
						assign rdata = rdata_r;
					end
				end
			end
			else begin : g_auto
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:245:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:248:13
								initial begin
									// Trace: src/VX_sp_ram.sv:248:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:250:13
								initial begin
									// Trace: src/VX_sp_ram.sv:251:17
									begin : sv2v_autoblock_13
										// Trace: src/VX_sp_ram.sv:251:22
										integer i;
										// Trace: src/VX_sp_ram.sv:251:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:252:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:257:21
						reg [ADDRW - 1:0] addr_r;
						// Trace: src/VX_sp_ram.sv:258:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:259:25
							if (read || write) begin
								// Trace: src/VX_sp_ram.sv:260:29
								if (write)
									// Trace: src/VX_sp_ram.sv:261:33
									begin : sv2v_autoblock_14
										// Trace: src/VX_sp_ram.sv:261:38
										integer i;
										// Trace: src/VX_sp_ram.sv:261:38
										for (i = 0; i < WRENW; i = i + 1)
											begin
												// Trace: src/VX_sp_ram.sv:262:33
												if (wren[i])
													// Trace: src/VX_sp_ram.sv:263:37
													ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
											end
									end
								// Trace: src/VX_sp_ram.sv:267:29
								addr_r <= addr;
							end
						// Trace: src/VX_sp_ram.sv:270:21
						assign rdata = ram[addr_r];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:272:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:275:13
								initial begin
									// Trace: src/VX_sp_ram.sv:275:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:277:13
								initial begin
									// Trace: src/VX_sp_ram.sv:278:17
									begin : sv2v_autoblock_15
										// Trace: src/VX_sp_ram.sv:278:22
										integer i;
										// Trace: src/VX_sp_ram.sv:278:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:279:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:284:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:285:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:286:25
							if (read || write) begin
								begin
									// Trace: src/VX_sp_ram.sv:287:29
									if (write) begin
										// Trace: src/VX_sp_ram.sv:288:33
										ram[addr] <= wdata;
										// Trace: src/VX_sp_ram.sv:289:33
										rdata_r <= wdata;
									end
									else
										// Trace: src/VX_sp_ram.sv:291:33
										rdata_r <= ram[addr];
								end
							end
						// Trace: src/VX_sp_ram.sv:295:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "R") begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:299:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:302:13
								initial begin
									// Trace: src/VX_sp_ram.sv:302:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:304:13
								initial begin
									// Trace: src/VX_sp_ram.sv:305:17
									begin : sv2v_autoblock_16
										// Trace: src/VX_sp_ram.sv:305:22
										integer i;
										// Trace: src/VX_sp_ram.sv:305:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:306:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:311:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:312:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:313:25
							if (read || write) begin
								// Trace: src/VX_sp_ram.sv:314:29
								if (write)
									// Trace: src/VX_sp_ram.sv:315:33
									begin : sv2v_autoblock_17
										// Trace: src/VX_sp_ram.sv:315:38
										integer i;
										// Trace: src/VX_sp_ram.sv:315:38
										for (i = 0; i < WRENW; i = i + 1)
											begin
												// Trace: src/VX_sp_ram.sv:316:33
												if (wren[i])
													// Trace: src/VX_sp_ram.sv:317:37
													ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
											end
									end
								// Trace: src/VX_sp_ram.sv:321:29
								rdata_r <= ram[addr];
							end
						// Trace: src/VX_sp_ram.sv:324:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:326:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:329:13
								initial begin
									// Trace: src/VX_sp_ram.sv:329:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:331:13
								initial begin
									// Trace: src/VX_sp_ram.sv:332:17
									begin : sv2v_autoblock_18
										// Trace: src/VX_sp_ram.sv:332:22
										integer i;
										// Trace: src/VX_sp_ram.sv:332:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:333:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:338:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:339:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:340:25
							if (read || write) begin
								// Trace: src/VX_sp_ram.sv:341:29
								if (write)
									// Trace: src/VX_sp_ram.sv:342:33
									ram[addr] <= wdata;
								// Trace: src/VX_sp_ram.sv:344:29
								rdata_r <= ram[addr];
							end
						// Trace: src/VX_sp_ram.sv:347:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "N") begin : g_no_change
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:351:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:354:13
								initial begin
									// Trace: src/VX_sp_ram.sv:354:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:356:13
								initial begin
									// Trace: src/VX_sp_ram.sv:357:17
									begin : sv2v_autoblock_19
										// Trace: src/VX_sp_ram.sv:357:22
										integer i;
										// Trace: src/VX_sp_ram.sv:357:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:358:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:363:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:364:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:365:25
							if (read || write) begin
								begin
									// Trace: src/VX_sp_ram.sv:366:29
									if (write)
										// Trace: src/VX_sp_ram.sv:367:33
										begin : sv2v_autoblock_20
											// Trace: src/VX_sp_ram.sv:367:38
											integer i;
											// Trace: src/VX_sp_ram.sv:367:38
											for (i = 0; i < WRENW; i = i + 1)
												begin
													// Trace: src/VX_sp_ram.sv:368:33
													if (wren[i])
														// Trace: src/VX_sp_ram.sv:369:37
														ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
												end
										end
									else
										// Trace: src/VX_sp_ram.sv:373:33
										rdata_r <= ram[addr];
								end
							end
						// Trace: src/VX_sp_ram.sv:377:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:379:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:382:13
								initial begin
									// Trace: src/VX_sp_ram.sv:382:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:384:13
								initial begin
									// Trace: src/VX_sp_ram.sv:385:17
									begin : sv2v_autoblock_21
										// Trace: src/VX_sp_ram.sv:385:22
										integer i;
										// Trace: src/VX_sp_ram.sv:385:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:386:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:391:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:392:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:393:25
							if (read || write) begin
								begin
									// Trace: src/VX_sp_ram.sv:394:29
									if (write)
										// Trace: src/VX_sp_ram.sv:395:33
										ram[addr] <= wdata;
									else
										// Trace: src/VX_sp_ram.sv:397:33
										rdata_r <= ram[addr];
								end
							end
						// Trace: src/VX_sp_ram.sv:401:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "U") begin : g_undefined
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:405:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:408:13
								initial begin
									// Trace: src/VX_sp_ram.sv:408:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:410:13
								initial begin
									// Trace: src/VX_sp_ram.sv:411:17
									begin : sv2v_autoblock_22
										// Trace: src/VX_sp_ram.sv:411:22
										integer i;
										// Trace: src/VX_sp_ram.sv:411:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:412:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:417:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:418:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:419:25
							if (write)
								// Trace: src/VX_sp_ram.sv:420:29
								begin : sv2v_autoblock_23
									// Trace: src/VX_sp_ram.sv:420:34
									integer i;
									// Trace: src/VX_sp_ram.sv:420:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:421:33
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:422:37
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_sp_ram.sv:427:29
								rdata_r <= ram[addr];
						end
						// Trace: src/VX_sp_ram.sv:430:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:432:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:435:13
								initial begin
									// Trace: src/VX_sp_ram.sv:435:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:437:13
								initial begin
									// Trace: src/VX_sp_ram.sv:438:17
									begin : sv2v_autoblock_24
										// Trace: src/VX_sp_ram.sv:438:22
										integer i;
										// Trace: src/VX_sp_ram.sv:438:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:439:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:444:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:445:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:446:25
							if (write)
								// Trace: src/VX_sp_ram.sv:447:29
								ram[addr] <= wdata;
							if (read)
								// Trace: src/VX_sp_ram.sv:450:29
								rdata_r <= ram[addr];
						end
						// Trace: src/VX_sp_ram.sv:453:21
						assign rdata = rdata_r;
					end
				end
			end
		end
		else begin : g_async
			if (FORCE_BRAM) begin : g_bram
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:461:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:464:13
								initial begin
									// Trace: src/VX_sp_ram.sv:464:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:466:13
								initial begin
									// Trace: src/VX_sp_ram.sv:467:17
									begin : sv2v_autoblock_25
										// Trace: src/VX_sp_ram.sv:467:22
										integer i;
										// Trace: src/VX_sp_ram.sv:467:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:468:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:473:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:474:25
							if (write)
								// Trace: src/VX_sp_ram.sv:475:29
								begin : sv2v_autoblock_26
									// Trace: src/VX_sp_ram.sv:475:34
									integer i;
									// Trace: src/VX_sp_ram.sv:475:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:476:33
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:477:37
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_sp_ram.sv:482:21
						assign rdata = ram[addr];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:484:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:487:13
								initial begin
									// Trace: src/VX_sp_ram.sv:487:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:489:13
								initial begin
									// Trace: src/VX_sp_ram.sv:490:17
									begin : sv2v_autoblock_27
										// Trace: src/VX_sp_ram.sv:490:22
										integer i;
										// Trace: src/VX_sp_ram.sv:490:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:491:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:496:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:497:25
							if (write)
								// Trace: src/VX_sp_ram.sv:498:29
								ram[addr] <= wdata;
						// Trace: src/VX_sp_ram.sv:501:21
						assign rdata = ram[addr];
					end
				end
				else begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:505:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:508:13
								initial begin
									// Trace: src/VX_sp_ram.sv:508:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:510:13
								initial begin
									// Trace: src/VX_sp_ram.sv:511:17
									begin : sv2v_autoblock_28
										// Trace: src/VX_sp_ram.sv:511:22
										integer i;
										// Trace: src/VX_sp_ram.sv:511:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:512:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:517:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:518:25
							if (write)
								// Trace: src/VX_sp_ram.sv:519:29
								begin : sv2v_autoblock_29
									// Trace: src/VX_sp_ram.sv:519:34
									integer i;
									// Trace: src/VX_sp_ram.sv:519:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:520:33
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:521:37
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_sp_ram.sv:526:21
						assign rdata = ram[addr];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:528:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:531:13
								initial begin
									// Trace: src/VX_sp_ram.sv:531:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:533:13
								initial begin
									// Trace: src/VX_sp_ram.sv:534:17
									begin : sv2v_autoblock_30
										// Trace: src/VX_sp_ram.sv:534:22
										integer i;
										// Trace: src/VX_sp_ram.sv:534:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:535:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:540:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:541:25
							if (write)
								// Trace: src/VX_sp_ram.sv:542:29
								ram[addr] <= wdata;
						// Trace: src/VX_sp_ram.sv:545:21
						assign rdata = ram[addr];
					end
				end
			end
			else begin : g_auto
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:551:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:554:13
								initial begin
									// Trace: src/VX_sp_ram.sv:554:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:556:13
								initial begin
									// Trace: src/VX_sp_ram.sv:557:17
									begin : sv2v_autoblock_31
										// Trace: src/VX_sp_ram.sv:557:22
										integer i;
										// Trace: src/VX_sp_ram.sv:557:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:558:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:563:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:564:25
							if (write)
								// Trace: src/VX_sp_ram.sv:565:29
								begin : sv2v_autoblock_32
									// Trace: src/VX_sp_ram.sv:565:34
									integer i;
									// Trace: src/VX_sp_ram.sv:565:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:566:33
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:567:37
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_sp_ram.sv:572:21
						assign rdata = ram[addr];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:574:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:577:13
								initial begin
									// Trace: src/VX_sp_ram.sv:577:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:579:13
								initial begin
									// Trace: src/VX_sp_ram.sv:580:17
									begin : sv2v_autoblock_33
										// Trace: src/VX_sp_ram.sv:580:22
										integer i;
										// Trace: src/VX_sp_ram.sv:580:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:581:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:586:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:587:25
							if (write)
								// Trace: src/VX_sp_ram.sv:588:29
								ram[addr] <= wdata;
						// Trace: src/VX_sp_ram.sv:591:21
						assign rdata = ram[addr];
					end
				end
				else begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:595:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:598:13
								initial begin
									// Trace: src/VX_sp_ram.sv:598:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:600:13
								initial begin
									// Trace: src/VX_sp_ram.sv:601:17
									begin : sv2v_autoblock_34
										// Trace: src/VX_sp_ram.sv:601:22
										integer i;
										// Trace: src/VX_sp_ram.sv:601:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:602:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:607:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:608:25
							if (write)
								// Trace: src/VX_sp_ram.sv:609:29
								begin : sv2v_autoblock_35
									// Trace: src/VX_sp_ram.sv:609:34
									integer i;
									// Trace: src/VX_sp_ram.sv:609:34
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:610:33
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:611:37
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_sp_ram.sv:616:21
						assign rdata = ram[addr];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:618:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:621:13
								initial begin
									// Trace: src/VX_sp_ram.sv:621:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:623:13
								initial begin
									// Trace: src/VX_sp_ram.sv:624:17
									begin : sv2v_autoblock_36
										// Trace: src/VX_sp_ram.sv:624:22
										integer i;
										// Trace: src/VX_sp_ram.sv:624:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:625:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:630:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:631:25
							if (write)
								// Trace: src/VX_sp_ram.sv:632:29
								ram[addr] <= wdata;
						// Trace: src/VX_sp_ram.sv:635:21
						assign rdata = ram[addr];
					end
				end
			end
		end
	endgenerate
endmodule
// removed module with interface ports: VX_operands
module fpnew_top_7C2B2_D4A54 (
	clk_i,
	rst_ni,
	operands_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	simd_mask_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:18:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	// removed localparam type fpnew_pkg_fpu_features_t
	localparam [42:0] fpnew_pkg_RV64D_Xsflt = 43'h000000207ff;
	parameter [42:0] Features = fpnew_pkg_RV64D_Xsflt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:19:13
	// removed localparam type fpnew_pkg_pipe_config_t
	// removed localparam type fpnew_pkg_unit_type_t
	localparam [31:0] fpnew_pkg_NUM_OPGROUPS = 4;
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unit_types_t
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unsigned_t
	// removed localparam type fpnew_pkg_fpu_implementation_t
	function automatic [159:0] sv2v_cast_B9240;
		input reg [159:0] inp;
		sv2v_cast_B9240 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 32) - 1:0] sv2v_cast_CDC93;
		input reg [((32'd4 * 32'd5) * 32) - 1:0] inp;
		sv2v_cast_CDC93 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 2) - 1:0] sv2v_cast_15FEF;
		input reg [((32'd4 * 32'd5) * 2) - 1:0] inp;
		sv2v_cast_15FEF = inp;
	endfunction
	localparam [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] fpnew_pkg_DEFAULT_NOREGS = {sv2v_cast_CDC93({fpnew_pkg_NUM_OPGROUPS {sv2v_cast_B9240(0)}}), sv2v_cast_15FEF({{fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}, {fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}}), 2'd0};
	parameter [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] Implementation = fpnew_pkg_DEFAULT_NOREGS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:21:13
	// removed localparam type fpnew_pkg_divsqrt_unit_t
	parameter [1:0] DivSqrtSel = 2'd2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:22:45
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:23:13
	parameter [31:0] TrueSIMDClass = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:24:13
	parameter [31:0] EnableSIMDMask = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:26:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:307:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:319:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:320:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:5
			begin : sv2v_autoblock_1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:323:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	function automatic signed [31:0] fpnew_pkg_minimum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:302:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:302:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:303:5
		fpnew_pkg_minimum = (a < b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_min_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:328:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:329:5
		reg [31:0] res;
		begin
			res = fpnew_pkg_max_fp_width(cfg);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:330:5
			begin : sv2v_autoblock_2
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:330:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:330:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:332:9
						res = $unsigned(fpnew_pkg_minimum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_min_fp_width = res;
		end
	endfunction
	function automatic [31:0] fpnew_pkg_max_num_lanes;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:405:49
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:405:69
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:405:86
		input reg vec;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:406:5
		fpnew_pkg_max_num_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg) : 1);
	endfunction
	localparam [31:0] NumLanes = fpnew_pkg_max_num_lanes(Features[42-:32], Features[8-:5], Features[10]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:27:27
	// removed localparam type MaskType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:28:14
	localparam [31:0] WIDTH = Features[42-:32];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:29:14
	localparam [31:0] NUM_OPERANDS = 3;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:31:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:32:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:34:3
	input wire [(NUM_OPERANDS * WIDTH) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:35:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:36:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:37:3
	input wire op_mod_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:38:3
	input wire [2:0] src_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:39:3
	input wire [2:0] dst_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:40:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:41:3
	input wire vectorial_op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:42:3
	input wire [TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:43:3
	input wire [NumLanes - 1:0] simd_mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:45:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:46:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:47:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:49:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:50:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:51:3
	output wire [TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:53:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:54:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:56:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:59:3
	localparam [31:0] NUM_OPGROUPS = fpnew_pkg_NUM_OPGROUPS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:60:3
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:65:3
	// removed localparam type output_t
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:72:3
	wire [3:0] opgrp_in_ready;
	wire [3:0] opgrp_out_valid;
	wire [3:0] opgrp_out_ready;
	wire [3:0] opgrp_ext;
	wire [3:0] opgrp_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:73:3
	wire [(4 * ((WIDTH + 5) + ((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)))) - 1:0] opgrp_outputs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:75:3
	wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:80:3
	// removed localparam type fpnew_pkg_opgroup_e
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [1:0] fpnew_pkg_get_opgroup;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:378:44
		input reg [3:0] op;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:379:5
		case (op)
			sv2v_cast_A53F3(0), sv2v_cast_A53F3(1), sv2v_cast_A53F3(2), sv2v_cast_A53F3(15), sv2v_cast_A53F3(3): fpnew_pkg_get_opgroup = 2'd0;
			sv2v_cast_A53F3(4), sv2v_cast_A53F3(5): fpnew_pkg_get_opgroup = 2'd1;
			sv2v_cast_A53F3(6), sv2v_cast_A53F3(7), sv2v_cast_A53F3(8), sv2v_cast_A53F3(9): fpnew_pkg_get_opgroup = 2'd2;
			sv2v_cast_A53F3(10), sv2v_cast_A53F3(11), sv2v_cast_A53F3(12), sv2v_cast_A53F3(13), sv2v_cast_A53F3(14): fpnew_pkg_get_opgroup = 2'd3;
			default: fpnew_pkg_get_opgroup = 2'd2;
		endcase
	endfunction
	assign in_ready_o = in_valid_i & opgrp_in_ready[fpnew_pkg_get_opgroup(op_i)];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:83:3
	genvar _gv_fmt_1;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_fmt_1 = 0; _gv_fmt_1 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_1 = _gv_fmt_1 + 1) begin : gen_nanbox_check
			localparam fmt = _gv_fmt_1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:84:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			if (Features[9] && (FP_WIDTH < WIDTH)) begin : check
				genvar _gv_op_1;
				for (_gv_op_1 = 0; _gv_op_1 < sv2v_cast_32_signed(NUM_OPERANDS); _gv_op_1 = _gv_op_1 + 1) begin : operands
					localparam op = _gv_op_1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:88:9
					assign is_boxed[(fmt * NUM_OPERANDS) + op] = (!vectorial_op_i ? operands_i[(op * WIDTH) + ((WIDTH - 1) >= FP_WIDTH ? WIDTH - 1 : ((WIDTH - 1) + ((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)) - 1)-:((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)] == {((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1) * 1 {1'sb1}} : 1'b1);
				end
			end
			else begin : no_check
				// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:93:7
				assign is_boxed[fmt * NUM_OPERANDS+:NUM_OPERANDS] = 1'sb1;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:98:3
	wire [NumLanes - 1:0] simd_mask;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:99:3
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	assign simd_mask = simd_mask_i | ~{NumLanes {sv2v_cast_1(EnableSIMDMask)}};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:104:3
	genvar _gv_opgrp_1;
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:389:48
		input reg [1:0] grp;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:390:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	generate
		for (_gv_opgrp_1 = 0; _gv_opgrp_1 < sv2v_cast_32_signed(NUM_OPGROUPS); _gv_opgrp_1 = _gv_opgrp_1 + 1) begin : gen_operation_groups
			localparam opgrp = _gv_opgrp_1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:105:5
			localparam [31:0] NUM_OPS = fpnew_pkg_num_operands(sv2v_cast_2(opgrp));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:106:5
			localparam [1:0] OpGroup = sv2v_cast_2(opgrp);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:107:5
			localparam [0:0] EnableVectors = Features[10];
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:108:5
			localparam [0:4] FpFmtMask = Features[8-:5];
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:109:5
			localparam [0:3] IntFmtMask = Features[3-:fpnew_pkg_NUM_INT_FORMATS];
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:110:5
			localparam [159:0] FmtPipeRegs = Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + (((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1)) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) - 1) - (32 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:160];
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:111:5
			localparam [9:0] FmtUnitTypes = Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) - 1) - (2 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:10];
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:112:5
			localparam [1:0] PipeConfig = Implementation[1-:2];
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:114:5
			wire in_valid;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:115:5
			reg [(NUM_FORMATS * NUM_OPS) - 1:0] input_boxed;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:117:5
			assign in_valid = in_valid_i & (fpnew_pkg_get_opgroup(op_i) == sv2v_cast_2(opgrp));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:120:5
			always @(*) begin : slice_inputs
				// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:121:7
				begin : sv2v_autoblock_3
					// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:121:12
					reg [31:0] fmt;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:121:12
					for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
						begin
							// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:122:9
							input_boxed[fmt * fpnew_pkg_num_operands(sv2v_cast_2(_gv_opgrp_1))+:fpnew_pkg_num_operands(sv2v_cast_2(_gv_opgrp_1))] = is_boxed[(fmt * NUM_OPERANDS) + (NUM_OPS - 1)-:NUM_OPS];
						end
				end
			end
			// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:125:5
			fpnew_opgroup_block_A87F3_05955 #(
				.TagType_TagType_TAG_WIDTH(TagType_TAG_WIDTH),
				.OpGroup(OpGroup),
				.Width(WIDTH),
				.EnableVectors(EnableVectors),
				.DivSqrtSel(DivSqrtSel),
				.FpFmtMask(FpFmtMask),
				.IntFmtMask(IntFmtMask),
				.FmtPipeRegs(FmtPipeRegs),
				.FmtUnitTypes(FmtUnitTypes),
				.PipeConfig(PipeConfig),
				.TrueSIMDClass(TrueSIMDClass)
			) i_opgroup_block(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i[WIDTH * ((NUM_OPS - 1) - (NUM_OPS - 1))+:WIDTH * NUM_OPS]),
				.is_boxed_i(input_boxed),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.simd_mask_i(simd_mask),
				.in_valid_i(in_valid),
				.in_ready_o(opgrp_in_ready[opgrp]),
				.flush_i(flush_i),
				.result_o(opgrp_outputs[(opgrp * ((WIDTH + 5) + ((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)))) + (WIDTH + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4))-:((WIDTH + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4)) >= (5 + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0)) ? ((WIDTH + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4)) - (5 + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((5 + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0)) - (WIDTH + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4))) + 1)]),
				.status_o(opgrp_outputs[(opgrp * ((WIDTH + 5) + ((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)))) + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4)-:((((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4) >= (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0) ? ((((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4) - (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0)) + 1 : ((((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0) - (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4)) + 1)]),
				.extension_bit_o(opgrp_ext[opgrp]),
				.tag_o(opgrp_outputs[(opgrp * ((WIDTH + 5) + ((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)))) + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) - 1)-:((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0))]),
				.out_valid_o(opgrp_out_valid[opgrp]),
				.out_ready_i(opgrp_out_ready[opgrp]),
				.busy_o(opgrp_busy[opgrp])
			);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:167:3
	wire [((WIDTH + 5) + ((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0))) - 1:0] arbiter_output;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:170:3
	localparam [31:0] sv2v_uu_i_arbiter_NumIn = NUM_OPGROUPS;
	localparam [31:0] sv2v_uu_i_arbiter_IdxWidth = $unsigned(2);
	// removed localparam type sv2v_uu_i_arbiter_rr_i
	localparam [sv2v_uu_i_arbiter_IdxWidth - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_CF21D_98F90 #(
		.DataType_TagType_TAG_WIDTH(TagType_TAG_WIDTH),
		.DataType_WIDTH(WIDTH),
		.NumIn(NUM_OPGROUPS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
		.req_i(opgrp_out_valid),
		.gnt_o(opgrp_out_ready),
		.data_i(opgrp_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:189:3
	assign result_o = arbiter_output[WIDTH + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4)-:((WIDTH + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4)) >= (5 + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0)) ? ((WIDTH + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4)) - (5 + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((5 + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0)) - (WIDTH + (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4))) + 1)];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:190:3
	assign status_o = arbiter_output[((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4-:((((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4) >= (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0) ? ((((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4) - (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0)) + 1 : ((((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 0) - (((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) + 4)) + 1)];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:191:3
	assign tag_o = arbiter_output[((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0)) - 1-:((TagType_TAG_WIDTH + 0) >= 0 ? TagType_TAG_WIDTH + 1 : 1 - (TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_top.sv:193:3
	assign busy_o = |opgrp_busy;
endmodule
module fpnew_opgroup_block_A87F3_05955 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	simd_mask_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:17:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:19:13
	parameter [31:0] Width = 32;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:20:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:21:13
	// removed localparam type fpnew_pkg_divsqrt_unit_t
	parameter [1:0] DivSqrtSel = 2'd2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:22:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtMask = 1'sb1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:23:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtMask = 1'sb1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:24:13
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	parameter [159:0] FmtPipeRegs = {fpnew_pkg_NUM_FP_FORMATS {32'd0}};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:25:13
	// removed localparam type fpnew_pkg_unit_type_t
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	parameter [9:0] FmtUnitTypes = {fpnew_pkg_NUM_FP_FORMATS {2'd1}};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:26:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:27:41
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:28:13
	parameter [31:0] TrueSIMDClass = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:30:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:31:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:389:48
		input reg [1:0] grp;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:390:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:32:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:307:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:319:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:320:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:5
			begin : sv2v_autoblock_1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:323:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	function automatic signed [31:0] fpnew_pkg_minimum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:302:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:302:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:303:5
		fpnew_pkg_minimum = (a < b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_min_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:328:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:329:5
		reg [31:0] res;
		begin
			res = fpnew_pkg_max_fp_width(cfg);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:330:5
			begin : sv2v_autoblock_2
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:330:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:330:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:332:9
						res = $unsigned(fpnew_pkg_minimum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_min_fp_width = res;
		end
	endfunction
	function automatic [31:0] fpnew_pkg_max_num_lanes;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:405:49
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:405:69
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:405:86
		input reg vec;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:406:5
		fpnew_pkg_max_num_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_max_num_lanes(Width, FpFmtMask, EnableVectors);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:33:27
	// removed localparam type MaskType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:35:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:36:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:38:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:39:3
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:40:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:41:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:42:3
	input wire op_mod_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:43:3
	input wire [2:0] src_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:44:3
	input wire [2:0] dst_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:45:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:46:3
	input wire vectorial_op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:47:3
	input wire [TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:48:3
	input wire [NUM_LANES - 1:0] simd_mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:50:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:51:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:52:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:54:3
	output wire [Width - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:55:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:56:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:57:3
	output wire [TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:59:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:60:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:62:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:68:3
	// removed localparam type output_t
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:76:3
	wire [4:0] fmt_in_ready;
	wire [4:0] fmt_out_valid;
	wire [4:0] fmt_out_ready;
	wire [4:0] fmt_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:77:3
	wire [(5 * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) - 1:0] fmt_outputs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:82:3
	assign in_ready_o = in_valid_i & fmt_in_ready[dst_fmt_i];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:87:3
	genvar _gv_fmt_2;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic fpnew_pkg_any_enabled_multi;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:476:46
		input reg [9:0] types;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:476:70
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:477:5
			begin : sv2v_autoblock_3
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:477:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:477:10
				begin : sv2v_autoblock_4
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_any_enabled_multi = 1'b1;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_any_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic [2:0] fpnew_pkg_get_first_enabled_multi;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:494:58
		input reg [9:0] types;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:494:82
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:495:5
			begin : sv2v_autoblock_5
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:495:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:495:10
				begin : sv2v_autoblock_6
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_get_first_enabled_multi = sv2v_cast_0BC43(i);
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_get_first_enabled_multi = sv2v_cast_0BC43(0);
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic fpnew_pkg_is_first_enabled_multi;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:484:51
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:485:51
		input reg [9:0] types;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:486:51
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:487:5
			begin : sv2v_autoblock_7
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:487:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:487:10
				begin : sv2v_autoblock_8
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:488:7
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_is_first_enabled_multi = sv2v_cast_0BC43(i) == fmt;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_is_first_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic [31:0] fpnew_pkg_num_lanes;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:400:45
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:400:65
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:400:82
		input reg vec;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:401:5
		fpnew_pkg_num_lanes = (vec ? width / fpnew_pkg_fp_width(fmt) : 1);
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	function automatic [((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) - 1:0] sv2v_cast_46BD0;
		input reg [((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) - 1:0] inp;
		sv2v_cast_46BD0 = inp;
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	generate
		for (_gv_fmt_2 = 0; _gv_fmt_2 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_2 = _gv_fmt_2 + 1) begin : gen_parallel_slices
			localparam fmt = _gv_fmt_2;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:89:5
			localparam [0:0] ANY_MERGED = fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:90:5
			localparam [0:0] IS_FIRST_MERGED = fpnew_pkg_is_first_enabled_multi(sv2v_cast_0BC43(fmt), FmtUnitTypes, FpFmtMask);
			if (FpFmtMask[fmt] && (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd1)) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:95:7
				localparam [2:0] FpFormat = sv2v_cast_0BC43(fmt);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:97:7
				wire in_valid;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:99:7
				assign in_valid = in_valid_i & (dst_fmt_i == fmt);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:102:7
				localparam [31:0] INTERNAL_LANES = fpnew_pkg_num_lanes(Width, sv2v_cast_0BC43(fmt), EnableVectors);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:103:7
				reg [INTERNAL_LANES - 1:0] mask_slice;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:104:7
				always @(*) begin : sv2v_autoblock_9
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:104:24
					reg signed [31:0] b;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:104:24
					for (b = 0; b < INTERNAL_LANES; b = b + 1)
						begin
							// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:104:60
							mask_slice[b] = simd_mask_i[(NUM_LANES / INTERNAL_LANES) * b];
						end
				end
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:106:7
				localparam [31:0] sv2v_uu_i_fmt_slice_NumPipeRegs = FmtPipeRegs[(4 - fmt) * 32+:32];
				localparam [31:0] sv2v_uu_i_fmt_slice_ExtRegEnaWidth = (sv2v_uu_i_fmt_slice_NumPipeRegs == 0 ? 1 : sv2v_uu_i_fmt_slice_NumPipeRegs);
				// removed localparam type sv2v_uu_i_fmt_slice_reg_ena_i
				localparam [sv2v_cast_32((sv2v_cast_32(FmtPipeRegs[(4 - _gv_fmt_2) * 32+:32]) == 0 ? 1 : sv2v_cast_32(FmtPipeRegs[(4 - _gv_fmt_2) * 32+:32]))) - 1:0] sv2v_uu_i_fmt_slice_ext_reg_ena_i_0 = 1'sb0;
				fpnew_opgroup_fmt_slice_F5668_FC739 #(
					.TagType_TagType_TagType_TAG_WIDTH(TagType_TagType_TAG_WIDTH),
					.OpGroup(OpGroup),
					.FpFormat(FpFormat),
					.Width(Width),
					.EnableVectors(EnableVectors),
					.NumPipeRegs(FmtPipeRegs[(4 - fmt) * 32+:32]),
					.PipeConfig(PipeConfig),
					.TrueSIMDClass(TrueSIMDClass)
				) i_fmt_slice(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.operands_i(operands_i),
					.is_boxed_i(is_boxed_i[fmt * NUM_OPERANDS+:NUM_OPERANDS]),
					.rnd_mode_i(rnd_mode_i),
					.op_i(op_i),
					.op_mod_i(op_mod_i),
					.vectorial_op_i(vectorial_op_i),
					.tag_i(tag_i),
					.simd_mask_i(mask_slice),
					.in_valid_i(in_valid),
					.in_ready_o(fmt_in_ready[fmt]),
					.flush_i(flush_i),
					.result_o(fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5))-:((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) >= (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) - (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5))) + 1)]),
					.status_o(fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)-:((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) >= (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) - (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) + 1)]),
					.extension_bit_o(fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)]),
					.tag_o(fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) - 1)-:((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0))]),
					.out_valid_o(fmt_out_valid[fmt]),
					.out_ready_i(fmt_out_ready[fmt]),
					.busy_o(fmt_busy[fmt]),
					.reg_ena_i(sv2v_uu_i_fmt_slice_ext_reg_ena_i_0)
				);
			end
			else if ((FpFmtMask[fmt] && ANY_MERGED) && !IS_FIRST_MERGED) begin : merged_unused
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:141:7
				localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:143:7
				assign fmt_in_ready[fmt] = fmt_in_ready[sv2v_cast_32_signed(FMT)];
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:145:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:146:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:148:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5))-:((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) >= (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) - (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5))) + 1)] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:149:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)-:((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) >= (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) - (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) + 1)] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:150:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)] = fpnew_pkg_DONT_CARE;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:151:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) - 1)-:((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0))] = sv2v_cast_46BD0(fpnew_pkg_DONT_CARE);
			end
			else if (!FpFmtMask[fmt] || (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd0)) begin : disable_fmt
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:155:7
				assign fmt_in_ready[fmt] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:156:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:157:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:159:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5))-:((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) >= (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) - (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5))) + 1)] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:160:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)-:((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) >= (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) - (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) + 1)] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:161:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)] = fpnew_pkg_DONT_CARE;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:162:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) - 1)-:((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0))] = sv2v_cast_46BD0(fpnew_pkg_DONT_CARE);
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:169:3
	function automatic [31:0] fpnew_pkg_get_num_regs_multi;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:502:54
		input reg [159:0] regs;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:503:54
		input reg [9:0] types;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:504:54
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:505:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:506:5
			begin : sv2v_autoblock_10
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:506:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:506:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:507:7
						if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2))
							// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:507:41
							res = fpnew_pkg_maximum(res, regs[(4 - i) * 32+:32]);
					end
			end
			fpnew_pkg_get_num_regs_multi = res;
		end
	endfunction
	generate
		if (fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask)) begin : gen_merged_slice
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:171:5
			localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:172:5
			localparam REG = fpnew_pkg_get_num_regs_multi(FmtPipeRegs, FmtUnitTypes, FpFmtMask);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:174:5
			wire in_valid;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:176:5
			assign in_valid = in_valid_i & (FmtUnitTypes[(4 - dst_fmt_i) * 2+:2] == 2'd2);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:178:5
			localparam [31:0] sv2v_uu_i_multifmt_slice_NumPipeRegs = REG;
			localparam [31:0] sv2v_uu_i_multifmt_slice_ExtRegEnaWidth = (sv2v_uu_i_multifmt_slice_NumPipeRegs == 0 ? 1 : sv2v_uu_i_multifmt_slice_NumPipeRegs);
			// removed localparam type sv2v_uu_i_multifmt_slice_reg_ena_i
			localparam [sv2v_uu_i_multifmt_slice_ExtRegEnaWidth - 1:0] sv2v_uu_i_multifmt_slice_ext_reg_ena_i_0 = 1'sb0;
			fpnew_opgroup_multifmt_slice_100B8_E15D3 #(
				.TagType_TagType_TagType_TAG_WIDTH(TagType_TagType_TAG_WIDTH),
				.OpGroup(OpGroup),
				.Width(Width),
				.FpFmtConfig(FpFmtMask),
				.IntFmtConfig(IntFmtMask),
				.EnableVectors(EnableVectors),
				.DivSqrtSel(DivSqrtSel),
				.NumPipeRegs(REG),
				.PipeConfig(PipeConfig)
			) i_multifmt_slice(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i),
				.is_boxed_i(is_boxed_i),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.simd_mask_i(simd_mask_i),
				.in_valid_i(in_valid),
				.in_ready_o(fmt_in_ready[FMT]),
				.flush_i(flush_i),
				.result_o(fmt_outputs[(FMT * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5))-:((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) >= (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) - (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5))) + 1)]),
				.status_o(fmt_outputs[(FMT * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)-:((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) >= (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) - (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) + 1)]),
				.extension_bit_o(fmt_outputs[(FMT * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)]),
				.tag_o(fmt_outputs[(FMT * ((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)))) + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) - 1)-:((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0))]),
				.out_valid_o(fmt_out_valid[FMT]),
				.out_ready_i(fmt_out_ready[FMT]),
				.busy_o(fmt_busy[FMT]),
				.reg_ena_i(sv2v_uu_i_multifmt_slice_ext_reg_ena_i_0)
			);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:220:3
	wire [((Width + 6) + ((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0))) - 1:0] arbiter_output;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:223:3
	localparam [31:0] sv2v_uu_i_arbiter_NumIn = NUM_FORMATS;
	localparam [31:0] sv2v_uu_i_arbiter_IdxWidth = $unsigned(3);
	// removed localparam type sv2v_uu_i_arbiter_rr_i
	localparam [sv2v_uu_i_arbiter_IdxWidth - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_4016C_91833 #(
		.DataType_TagType_TagType_TAG_WIDTH(TagType_TagType_TAG_WIDTH),
		.DataType_Width(Width),
		.NumIn(NUM_FORMATS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
		.req_i(fmt_out_valid),
		.gnt_o(fmt_out_ready),
		.data_i(fmt_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:242:3
	assign result_o = arbiter_output[Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)-:((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) >= (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) - (6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((6 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (Width + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5))) + 1)];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:243:3
	assign status_o = arbiter_output[((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5-:((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) >= (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) ? ((((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5) - (1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0))) + 1 : ((1 + (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0)) - (((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 5)) + 1)];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:244:3
	assign extension_bit_o = arbiter_output[((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) + 0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:245:3
	assign tag_o = arbiter_output[((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0)) - 1-:((TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_block.sv:247:3
	assign busy_o = |fmt_busy;
endmodule
module fpnew_opgroup_multifmt_slice_100B8_E15D3 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	simd_mask_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o,
	reg_ena_i
);
	// removed localparam type TagType_TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:19:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd3;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:20:13
	parameter [31:0] Width = 64;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:22:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:23:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtConfig = 1'sb1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:24:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:25:13
	// removed localparam type fpnew_pkg_divsqrt_unit_t
	parameter [1:0] DivSqrtSel = 2'd2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:26:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:27:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:28:13
	parameter [0:0] ExtRegEna = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:29:39
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:31:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:389:48
		input reg [1:0] grp;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:390:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:32:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:33:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:307:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:319:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:320:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:5
			begin : sv2v_autoblock_1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:323:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	function automatic signed [31:0] fpnew_pkg_minimum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:302:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:302:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:303:5
		fpnew_pkg_minimum = (a < b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_min_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:328:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:329:5
		reg [31:0] res;
		begin
			res = fpnew_pkg_max_fp_width(cfg);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:330:5
			begin : sv2v_autoblock_2
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:330:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:330:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:332:9
						res = $unsigned(fpnew_pkg_minimum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_min_fp_width = res;
		end
	endfunction
	function automatic [31:0] fpnew_pkg_max_num_lanes;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:405:49
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:405:69
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:405:86
		input reg vec;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:406:5
		fpnew_pkg_max_num_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg) : 1);
	endfunction
	localparam [31:0] NUM_SIMD_LANES = fpnew_pkg_max_num_lanes(Width, FpFmtConfig, EnableVectors);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:34:27
	// removed localparam type MaskType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:35:14
	localparam [31:0] ExtRegEnaWidth = (NumPipeRegs == 0 ? 1 : NumPipeRegs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:37:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:38:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:40:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:41:3
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:42:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:43:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:44:3
	input wire op_mod_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:45:3
	input wire [2:0] src_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:46:3
	input wire [2:0] dst_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:47:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:48:3
	input wire vectorial_op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:49:3
	input wire [TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:50:3
	input wire [NUM_SIMD_LANES - 1:0] simd_mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:52:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:53:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:54:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:56:3
	output wire [Width - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:57:3
	// removed localparam type fpnew_pkg_status_t
	output reg [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:58:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:59:3
	output wire [TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:61:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:62:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:64:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:66:3
	input wire [ExtRegEnaWidth - 1:0] reg_ena_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:69:3
	generate
		if (OpGroup == 2'd1) begin : genblk1
			if ((DivSqrtSel == 2'd1) && !((FpFmtConfig[0] == 1) && (FpFmtConfig[1:4] == {4 {1'sb0}}))) begin : genblk1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:71:7
				$fatal(1, "T-Head-based DivSqrt unit supported only in FP32-only configurations. Set DivSqrtSel = THMULTI or DivSqrtSel = PULP to use a multi-format divider");
			end
			else if ((DivSqrtSel == 2'd2) && (FpFmtConfig[3] == 1'b1)) begin : genblk1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:74:7
				$warning("The DivSqrt unit of C910 (instantiated by DivSqrtSel = THMULTI) does not support FP8. Please use the PULP DivSqrt unit when in need of div/sqrt operations on FP8.");
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:79:3
	localparam [31:0] MAX_FP_WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:80:3
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:88:45
		input reg [1:0] ifmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:89:5
		case (ifmt)
			sv2v_cast_87CC5(0): fpnew_pkg_int_width = 8;
			sv2v_cast_87CC5(1): fpnew_pkg_int_width = 16;
			sv2v_cast_87CC5(2): fpnew_pkg_int_width = 32;
			sv2v_cast_87CC5(3): fpnew_pkg_int_width = 64;
			default: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:96:9
				$fatal(1, "Invalid INT format supplied");
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:100:9
				fpnew_pkg_int_width = sv2v_cast_87CC5(0);
			end
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:366:49
		input reg [0:3] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:367:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:368:5
			begin : sv2v_autoblock_3
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:368:10
				reg signed [31:0] ifmt;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:368:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:369:7
						if (cfg[ifmt])
							// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:369:22
							res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)));
					end
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:81:3
	localparam [31:0] NUM_LANES = fpnew_pkg_max_num_lanes(Width, FpFmtConfig, 1'b1);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:82:3
	function automatic [31:0] fpnew_pkg_num_divsqrt_lanes;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:410:53
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:410:73
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:410:90
		input reg vec;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:410:101
		input reg [1:0] DivSqrtSel;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:411:5
		reg [0:4] cfg_tmp;
		begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:412:5
			cfg_tmp = (DivSqrtSel == 2'd2 ? cfg & 5'b11101 : cfg);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:413:5
			fpnew_pkg_num_divsqrt_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg_tmp) : 1);
		end
	endfunction
	localparam [31:0] NUM_DIVSQRT_LANES = fpnew_pkg_num_divsqrt_lanes(Width, FpFmtConfig, 1'b1, DivSqrtSel);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:83:3
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:85:3
	localparam [31:0] FMT_BITS = fpnew_pkg_maximum(3, 2);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:87:3
	localparam [31:0] AUX_BITS = FMT_BITS + 2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:89:3
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	wire [NUM_LANES - 1:0] divsqrt_done;
	wire [NUM_LANES - 1:0] divsqrt_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:90:3
	wire vectorial_op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:91:3
	wire [FMT_BITS - 1:0] dst_fmt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:92:3
	wire [AUX_BITS - 1:0] aux_data;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:95:3
	wire dst_fmt_is_int;
	wire dst_is_cpk;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:96:3
	wire [1:0] dst_vec_op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:97:3
	wire [2:0] target_aux_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:98:3
	wire is_up_cast;
	wire is_down_cast;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:100:3
	wire [(NUM_FORMATS * Width) - 1:0] fmt_slice_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:101:3
	wire [(NUM_INT_FORMATS * Width) - 1:0] ifmt_slice_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:103:3
	wire [Width - 1:0] conv_target_d;
	wire [Width - 1:0] conv_target_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:105:3
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:106:3
	wire [NUM_LANES - 1:0] lane_ext_bit;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:107:3
	wire [((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? (NUM_LANES * (TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : (NUM_LANES * (1 - (TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TAG_WIDTH - 1)):((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0)] lane_tags;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:108:3
	wire [NUM_LANES - 1:0] lane_masks;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:109:3
	wire [(NUM_LANES * AUX_BITS) - 1:0] lane_aux;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:110:3
	wire [NUM_LANES - 1:0] lane_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:112:3
	wire result_is_vector;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:113:3
	wire [FMT_BITS - 1:0] result_fmt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:114:3
	wire result_fmt_is_int;
	wire result_is_cpk;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:115:3
	wire [1:0] result_vec_op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:117:3
	wire simd_synch_rdy;
	wire simd_synch_done;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:122:3
	assign in_ready_o = lane_in_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:123:3
	assign vectorial_op = vectorial_op_i & EnableVectors;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:126:3
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	assign dst_fmt_is_int = (OpGroup == 2'd3) & (op_i == sv2v_cast_A53F3(11));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:127:3
	assign dst_is_cpk = (OpGroup == 2'd3) & ((op_i == sv2v_cast_A53F3(13)) || (op_i == sv2v_cast_A53F3(14)));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:129:3
	assign dst_vec_op = (OpGroup == 2'd3) & {op_i == sv2v_cast_A53F3(14), op_mod_i};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:131:3
	assign is_up_cast = fpnew_pkg_fp_width(dst_fmt_i) > fpnew_pkg_fp_width(src_fmt_i);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:132:3
	assign is_down_cast = fpnew_pkg_fp_width(dst_fmt_i) < fpnew_pkg_fp_width(src_fmt_i);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:135:3
	assign dst_fmt = (dst_fmt_is_int ? int_fmt_i : dst_fmt_i);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:138:3
	assign aux_data = {dst_fmt_is_int, vectorial_op, dst_fmt};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:139:3
	assign target_aux_d = {dst_vec_op, dst_is_cpk};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:142:3
	generate
		if (OpGroup == 2'd3) begin : conv_target
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:143:5
			assign conv_target_d = (dst_is_cpk ? operands_i[2 * Width+:Width] : operands_i[Width+:Width]);
		end
		else begin : not_conv_target
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:145:5
			assign conv_target_d = 1'sb0;
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:149:3
	reg [4:0] is_boxed_1op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:150:3
	reg [9:0] is_boxed_2op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:152:3
	always @(*) begin : boxed_2op
		// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:153:5
		begin : sv2v_autoblock_4
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:153:10
			reg signed [31:0] fmt;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:153:10
			for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
				begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:154:7
					is_boxed_1op[fmt] = is_boxed_i[fmt * NUM_OPERANDS];
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:155:7
					is_boxed_2op[fmt * 2+:2] = is_boxed_i[(fmt * NUM_OPERANDS) + 1-:2];
				end
		end
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:162:3
	genvar _gv_lane_1;
	localparam [0:4] fpnew_pkg_CPK_FORMATS = 5'b11000;
	function automatic [0:4] fpnew_pkg_get_conv_lane_formats;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:446:56
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:447:56
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:448:56
		input reg [31:0] lane_no;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:449:5
		reg [0:4] res;
		begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:450:5
			begin : sv2v_autoblock_5
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:450:10
				reg [31:0] fmt;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:450:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:452:7
						res[fmt] = cfg[fmt] && (((width / fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))) > lane_no) || (fpnew_pkg_CPK_FORMATS[fmt] && (lane_no < 2)));
					end
			end
			fpnew_pkg_get_conv_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_conv_lane_int_formats;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:458:61
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:459:61
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:460:61
		input reg [0:3] icfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:461:61
		input reg [31:0] lane_no;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:462:5
		reg [0:3] res;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:463:5
		reg [0:4] lanefmts;
		begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:464:5
			res = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:465:5
			lanefmts = fpnew_pkg_get_conv_lane_formats(width, cfg, lane_no);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:467:5
			begin : sv2v_autoblock_6
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:467:10
				reg [31:0] ifmt;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:467:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_7
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:468:12
						reg [31:0] fmt;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:468:12
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							begin
								// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:470:9
								res[ifmt] = res[ifmt] | ((icfg[ifmt] && lanefmts[fmt]) && (fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt)) == fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt))));
							end
					end
			end
			fpnew_pkg_get_conv_lane_int_formats = res;
		end
	endfunction
	function automatic [0:4] fpnew_pkg_get_lane_formats;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:417:51
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:418:51
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:419:51
		input reg [31:0] lane_no;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:420:5
		reg [0:4] res;
		begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:421:5
			begin : sv2v_autoblock_8
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:421:10
				reg [31:0] fmt;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:421:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:423:7
						res[fmt] = cfg[fmt] & ((width / fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))) > lane_no);
					end
			end
			fpnew_pkg_get_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_lane_int_formats;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:428:56
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:429:56
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:430:56
		input reg [0:3] icfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:431:56
		input reg [31:0] lane_no;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:432:5
		reg [0:3] res;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:433:5
		reg [0:4] lanefmts;
		begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:434:5
			res = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:435:5
			lanefmts = fpnew_pkg_get_lane_formats(width, cfg, lane_no);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:437:5
			begin : sv2v_autoblock_9
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:437:10
				reg [31:0] ifmt;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:437:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_10
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:438:12
						reg [31:0] fmt;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:438:12
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							if (fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt)) == fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)))
								// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:441:11
								res[ifmt] = res[ifmt] | (icfg[ifmt] && lanefmts[fmt]);
					end
			end
			fpnew_pkg_get_lane_int_formats = res;
		end
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [4:0] sv2v_cast_F8FCA;
		input reg [4:0] inp;
		sv2v_cast_F8FCA = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_lane_1 = 0; _gv_lane_1 < sv2v_cast_32_signed(NUM_LANES); _gv_lane_1 = _gv_lane_1 + 1) begin : gen_num_lanes
			localparam lane = _gv_lane_1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:163:5
			localparam [31:0] LANE = $unsigned(lane);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:165:5
			localparam [0:4] ACTIVE_FORMATS = fpnew_pkg_get_lane_formats(Width, FpFmtConfig, LANE);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:167:5
			localparam [0:3] ACTIVE_INT_FORMATS = fpnew_pkg_get_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:169:5
			localparam [31:0] MAX_WIDTH = fpnew_pkg_max_fp_width(ACTIVE_FORMATS);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:172:5
			localparam [0:4] CONV_FORMATS = fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, LANE);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:174:5
			localparam [0:3] CONV_INT_FORMATS = fpnew_pkg_get_conv_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:176:5
			localparam [31:0] CONV_WIDTH = fpnew_pkg_max_fp_width(CONV_FORMATS);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:179:5
			localparam [0:4] LANE_FORMATS = (OpGroup == 2'd3 ? CONV_FORMATS : ACTIVE_FORMATS);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:181:5
			localparam [31:0] LANE_WIDTH = (OpGroup == 2'd3 ? CONV_WIDTH : MAX_WIDTH);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:183:5
			wire [LANE_WIDTH - 1:0] local_result;
			if ((lane == 0) || (EnableVectors & !((OpGroup == 2'd1) && (lane >= NUM_DIVSQRT_LANES)))) begin : active_lane
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:187:7
				wire in_valid;
				wire out_valid;
				wire out_ready;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:189:7
				reg [(NUM_OPERANDS * LANE_WIDTH) - 1:0] local_operands;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:190:7
				wire [LANE_WIDTH - 1:0] op_result;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:191:7
				wire [4:0] op_status;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:193:7
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:196:7
				always @(*) begin : prepare_input
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:197:9
					begin : sv2v_autoblock_11
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:197:14
						reg [31:0] i;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:197:14
						for (i = 0; i < NUM_OPERANDS; i = i + 1)
							begin
								// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:198:11
								if (i == 2)
									// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:199:13
									local_operands[i * (OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))))+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))))] = operands_i[i * Width+:Width] >> (LANE * fpnew_pkg_fp_width((op_i == sv2v_cast_A53F3(15) ? src_fmt_i : dst_fmt_i)));
								else
									// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:201:13
									local_operands[i * (OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))))+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))))] = operands_i[i * Width+:Width] >> (LANE * fpnew_pkg_fp_width(src_fmt_i));
							end
					end
					if (OpGroup == 2'd3) begin
						begin
							// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:208:11
							if (op_i == sv2v_cast_A53F3(12))
								// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:209:13
								local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))))] = operands_i[0+:Width] >> (LANE * fpnew_pkg_int_width(int_fmt_i));
							else if (op_i == sv2v_cast_A53F3(10)) begin
								begin
									// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:212:13
									if ((vectorial_op && op_mod_i) && is_up_cast)
										// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:213:15
										local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))))] = operands_i[0+:Width] >> ((LANE * fpnew_pkg_fp_width(src_fmt_i)) + (MAX_FP_WIDTH / 2));
								end
							end
							else if (dst_is_cpk) begin
								begin
									// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:218:13
									if (lane == 1)
										// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:219:15
										local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))))] = operands_i[Width + (LANE_WIDTH - 1)-:LANE_WIDTH];
								end
							end
						end
					end
				end
				if (OpGroup == 2'd0) begin : lane_instance
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:227:9
					fpnew_fma_multi_6D055_6E71C #(
						.AuxType_AUX_BITS(AUX_BITS),
						.TagType_TagType_TagType_TagType_TAG_WIDTH(TagType_TagType_TagType_TAG_WIDTH),
						.FpFmtConfig(LANE_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_fma_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.src2_fmt_i((op_i == sv2v_cast_A53F3(15) ? src_fmt_i : dst_fmt_i)),
						.dst_fmt_i(dst_fmt_i),
						.tag_i(tag_i),
						.mask_i(simd_mask_i[lane]),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + (lane * ((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))]),
						.mask_o(lane_masks[lane]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane]),
						.reg_ena_i(reg_ena_i)
					);
				end
				else if (OpGroup == 2'd1) begin : lane_instance
					if (((DivSqrtSel == 2'd1) && LANE_FORMATS[0]) && (LANE_FORMATS[1:4] == {4 {1'sb0}})) begin : gen_th32_e906_divsqrt
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:265:11
						fpnew_divsqrt_th_32_2BDD9_C9EC9 #(
							.AuxType_AUX_BITS(AUX_BITS),
							.TagType_TagType_TagType_TagType_TAG_WIDTH(TagType_TagType_TagType_TAG_WIDTH),
							.NumPipeRegs(NumPipeRegs),
							.PipeConfig(PipeConfig)
						) i_fpnew_divsqrt_multi_th(
							.clk_i(clk_i),
							.rst_ni(rst_ni),
							.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1))))) * 2]),
							.is_boxed_i(is_boxed_2op),
							.rnd_mode_i(rnd_mode_i),
							.op_i(op_i),
							.tag_i(tag_i),
							.mask_i(simd_mask_i[lane]),
							.aux_i(aux_data),
							.in_valid_i(in_valid),
							.in_ready_o(lane_in_ready[lane]),
							.flush_i(flush_i),
							.result_o(op_result),
							.status_o(op_status),
							.extension_bit_o(lane_ext_bit[lane]),
							.tag_o(lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + (lane * ((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))]),
							.mask_o(lane_masks[lane]),
							.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
							.out_valid_o(out_valid),
							.out_ready_i(out_ready),
							.busy_o(lane_busy[lane]),
							.reg_ena_i(reg_ena_i)
						);
					end
					else if (DivSqrtSel == 2'd2) begin : gen_thmulti_c910_divsqrt
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:295:11
						fpnew_divsqrt_th_64_multi_5F898_8E3CD #(
							.AuxType_AUX_BITS(AUX_BITS),
							.TagType_TagType_TagType_TagType_TAG_WIDTH(TagType_TagType_TagType_TAG_WIDTH),
							.FpFmtConfig(LANE_FORMATS),
							.NumPipeRegs(NumPipeRegs),
							.PipeConfig(PipeConfig)
						) i_fpnew_divsqrt_th_64_c910(
							.clk_i(clk_i),
							.rst_ni(rst_ni),
							.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1))))) * 2]),
							.is_boxed_i(is_boxed_2op),
							.rnd_mode_i(rnd_mode_i),
							.op_i(op_i),
							.dst_fmt_i(dst_fmt_i),
							.tag_i(tag_i),
							.mask_i(simd_mask_i[lane]),
							.aux_i(aux_data),
							.vectorial_op_i(vectorial_op),
							.in_valid_i(in_valid),
							.in_ready_o(lane_in_ready[lane]),
							.divsqrt_done_o(divsqrt_done[lane]),
							.simd_synch_done_i(simd_synch_done),
							.divsqrt_ready_o(divsqrt_ready[lane]),
							.simd_synch_rdy_i(simd_synch_rdy),
							.flush_i(flush_i),
							.result_o(op_result),
							.status_o(op_status),
							.extension_bit_o(lane_ext_bit[lane]),
							.tag_o(lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + (lane * ((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))]),
							.mask_o(lane_masks[lane]),
							.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
							.out_valid_o(out_valid),
							.out_ready_i(out_ready),
							.busy_o(lane_busy[lane]),
							.reg_ena_i(reg_ena_i)
						);
					end
					else begin : gen_pulp_divsqrt
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:332:11
						fpnew_divsqrt_multi_68C3A_AC02A #(
							.AuxType_AUX_BITS(AUX_BITS),
							.TagType_TagType_TagType_TagType_TAG_WIDTH(TagType_TagType_TagType_TAG_WIDTH),
							.FpFmtConfig(LANE_FORMATS),
							.NumPipeRegs(NumPipeRegs),
							.PipeConfig(PipeConfig)
						) i_fpnew_divsqrt_multi(
							.clk_i(clk_i),
							.rst_ni(rst_ni),
							.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1))))) * 2]),
							.is_boxed_i(is_boxed_2op),
							.rnd_mode_i(rnd_mode_i),
							.op_i(op_i),
							.dst_fmt_i(dst_fmt_i),
							.tag_i(tag_i),
							.mask_i(simd_mask_i[lane]),
							.aux_i(aux_data),
							.vectorial_op_i(vectorial_op),
							.in_valid_i(in_valid),
							.in_ready_o(lane_in_ready[lane]),
							.divsqrt_done_o(divsqrt_done[lane]),
							.simd_synch_done_i(simd_synch_done),
							.divsqrt_ready_o(divsqrt_ready[lane]),
							.simd_synch_rdy_i(simd_synch_rdy),
							.flush_i(flush_i),
							.result_o(op_result),
							.status_o(op_status),
							.extension_bit_o(lane_ext_bit[lane]),
							.tag_o(lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + (lane * ((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))]),
							.mask_o(lane_masks[lane]),
							.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
							.out_valid_o(out_valid),
							.out_ready_i(out_ready),
							.busy_o(lane_busy[lane]),
							.reg_ena_i(reg_ena_i)
						);
					end
				end
				else if (OpGroup == 2'd2) begin
					;
				end
				else if (OpGroup == 2'd3) begin : lane_instance
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:372:9
					fpnew_cast_multi_ACFE7_57164 #(
						.AuxType_AUX_BITS(AUX_BITS),
						.TagType_TagType_TagType_TagType_TAG_WIDTH(TagType_TagType_TagType_TAG_WIDTH),
						.FpFmtConfig(LANE_FORMATS),
						.IntFmtConfig(CONV_INT_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_cast_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))))]),
						.is_boxed_i(is_boxed_1op),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.dst_fmt_i(dst_fmt_i),
						.int_fmt_i(int_fmt_i),
						.tag_i(tag_i),
						.mask_i(simd_mask_i[lane]),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + (lane * ((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))]),
						.mask_o(lane_masks[lane]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane]),
						.reg_ena_i(reg_ena_i)
					);
				end
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:410:7
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:411:7
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:414:7
				assign local_result = (lane_out_valid[lane] | ExtRegEna ? op_result : {(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1))))) : fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(_gv_lane_1)))))) {lane_ext_bit[0]}});
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:415:7
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] | ExtRegEna ? op_status : {5 {1'sb0}});
			end
			else begin : inactive_lane
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:419:7
				assign lane_out_valid[lane] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:420:7
				assign lane_in_ready[lane] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:421:7
				assign lane_aux[lane * AUX_BITS+:AUX_BITS] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:422:7
				assign lane_masks[lane] = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:423:7
				assign lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + (lane * ((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:424:7
				assign divsqrt_done[lane] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:425:7
				assign divsqrt_ready[lane] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:426:7
				assign lane_ext_bit[lane] = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:427:7
				assign local_result = {LANE_WIDTH {lane_ext_bit[0]}};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:428:7
				assign lane_status[lane * 5+:5] = 1'sb0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:429:7
				assign lane_busy[lane] = 1'b0;
			end
			genvar _gv_fmt_3;
			for (_gv_fmt_3 = 0; _gv_fmt_3 < NUM_FORMATS; _gv_fmt_3 = _gv_fmt_3 + 1) begin : pack_fp_result
				localparam fmt = _gv_fmt_3;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:435:7
				localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
				if (ACTIVE_FORMATS[fmt]) begin : genblk1
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:438:9
					assign fmt_slice_result[(fmt * Width) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((LANE + 1) * FP_WIDTH) - 1 : ((((LANE + 1) * FP_WIDTH) - 1) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)] = local_result[FP_WIDTH - 1:0];
				end
				else if (((LANE + 1) * FP_WIDTH) <= Width) begin : genblk1
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:441:9
					assign fmt_slice_result[(fmt * Width) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((LANE + 1) * FP_WIDTH) - 1 : ((((LANE + 1) * FP_WIDTH) - 1) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)] = {((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1) {lane_ext_bit[LANE]}};
				end
				else if ((LANE * FP_WIDTH) < Width) begin : genblk1
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:444:9
					assign fmt_slice_result[(fmt * Width) + ((Width - 1) >= (LANE * FP_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1)] = {((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1) {lane_ext_bit[LANE]}};
				end
			end
			if (OpGroup == 2'd3) begin : int_results_enabled
				genvar _gv_ifmt_1;
				for (_gv_ifmt_1 = 0; _gv_ifmt_1 < NUM_INT_FORMATS; _gv_ifmt_1 = _gv_ifmt_1 + 1) begin : pack_int_result
					localparam ifmt = _gv_ifmt_1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:453:9
					localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
					if (ACTIVE_INT_FORMATS[ifmt]) begin : genblk1
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:455:11
						assign ifmt_slice_result[(ifmt * Width) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((LANE + 1) * INT_WIDTH) - 1 : ((((LANE + 1) * INT_WIDTH) - 1) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)] = local_result[INT_WIDTH - 1:0];
					end
					else if (((LANE + 1) * INT_WIDTH) <= Width) begin : genblk1
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:458:11
						assign ifmt_slice_result[(ifmt * Width) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((LANE + 1) * INT_WIDTH) - 1 : ((((LANE + 1) * INT_WIDTH) - 1) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)] = 1'sb0;
					end
					else if ((LANE * INT_WIDTH) < Width) begin : genblk1
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:460:11
						assign ifmt_slice_result[(ifmt * Width) + ((Width - 1) >= (LANE * INT_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (LANE * INT_WIDTH) ? ((Width - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (LANE * INT_WIDTH) ? ((Width - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (Width - 1)) + 1)] = 1'sb0;
					end
				end
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:467:3
	genvar _gv_fmt_4;
	generate
		for (_gv_fmt_4 = 0; _gv_fmt_4 < NUM_FORMATS; _gv_fmt_4 = _gv_fmt_4 + 1) begin : extend_fp_result
			localparam fmt = _gv_fmt_4;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:469:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			if ((NUM_LANES * FP_WIDTH) < Width) begin : genblk1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:471:7
				assign fmt_slice_result[(fmt * Width) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)] = {((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1) {lane_ext_bit[0]}};
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:474:3
	genvar _gv_ifmt_2;
	generate
		for (_gv_ifmt_2 = 0; _gv_ifmt_2 < NUM_INT_FORMATS; _gv_ifmt_2 = _gv_ifmt_2 + 1) begin : extend_or_mute_int_result
			localparam ifmt = _gv_ifmt_2;
			if (OpGroup != 2'd3) begin : mute_int_result
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:477:7
				assign ifmt_slice_result[ifmt * Width+:Width] = 1'sb0;
			end
			else begin : extend_int_result
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:482:7
				localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
				if ((NUM_LANES * INT_WIDTH) < Width) begin : genblk1
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:484:9
					assign ifmt_slice_result[(ifmt * Width) + ((Width - 1) >= (NUM_LANES * INT_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (NUM_LANES * INT_WIDTH) ? ((Width - 1) - (NUM_LANES * INT_WIDTH)) + 1 : ((NUM_LANES * INT_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (NUM_LANES * INT_WIDTH) ? ((Width - 1) - (NUM_LANES * INT_WIDTH)) + 1 : ((NUM_LANES * INT_WIDTH) - (Width - 1)) + 1)] = 1'sb0;
				end
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:489:3
	generate
		if (OpGroup == 2'd3) begin : target_regs
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:491:5
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * Width) + ((NumPipeRegs * Width) - 1) : ((NumPipeRegs + 1) * Width) - 1):(0 >= NumPipeRegs ? NumPipeRegs * Width : 0)] byp_pipe_target_q;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:492:5
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * 3) + ((NumPipeRegs * 3) - 1) : ((NumPipeRegs + 1) * 3) - 1):(0 >= NumPipeRegs ? NumPipeRegs * 3 : 0)] byp_pipe_aux_q;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:493:5
			reg [0:NumPipeRegs] byp_pipe_valid_q;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:495:5
			wire [0:NumPipeRegs] byp_pipe_ready;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:498:5
			wire [Width * 1:1] sv2v_tmp_FBD8C;
			assign sv2v_tmp_FBD8C = conv_target_d;
			always @(*) byp_pipe_target_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * Width+:Width] = sv2v_tmp_FBD8C;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:499:5
			wire [3:1] sv2v_tmp_A0A5D;
			assign sv2v_tmp_A0A5D = target_aux_d;
			always @(*) byp_pipe_aux_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * 3+:3] = sv2v_tmp_A0A5D;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:500:5
			wire [1:1] sv2v_tmp_49222;
			assign sv2v_tmp_49222 = in_valid_i & vectorial_op;
			always @(*) byp_pipe_valid_q[0] = sv2v_tmp_49222;
			genvar _gv_i_218;
			for (_gv_i_218 = 0; _gv_i_218 < NumPipeRegs; _gv_i_218 = _gv_i_218 + 1) begin : gen_bypass_pipeline
				localparam i = _gv_i_218;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:504:7
				wire reg_ena;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:508:7
				assign byp_pipe_ready[i] = byp_pipe_ready[i + 1] | ~byp_pipe_valid_q[i + 1];
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:510:254
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:510:332
					if (!rst_ni)
						// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:510:410
						byp_pipe_valid_q[i + 1] <= 1'b0;
					else
						// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:510:562
						byp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (byp_pipe_ready[i] ? byp_pipe_valid_q[i] : byp_pipe_valid_q[i + 1]));
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:512:7
				assign reg_ena = (byp_pipe_ready[i] & byp_pipe_valid_q[i]) | reg_ena_i[i];
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:514:71
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:514:127
					if (!rst_ni)
						// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:514:183
						byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= 1'sb0;
					else
						// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:514:291
						byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= (reg_ena ? byp_pipe_target_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * Width+:Width] : byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width]);
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:515:71
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:515:127
					if (!rst_ni)
						// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:515:183
						byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= 1'sb0;
					else
						// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:515:291
						byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= (reg_ena ? byp_pipe_aux_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * 3+:3] : byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3]);
			end
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:518:5
			assign byp_pipe_ready[NumPipeRegs] = out_ready_i & result_is_vector;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:520:5
			assign conv_target_q = byp_pipe_target_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * Width+:Width];
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:523:5
			assign {result_vec_op, result_is_cpk} = byp_pipe_aux_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * 3+:3];
		end
		else begin : no_conv
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:525:5
			assign {result_vec_op, result_is_cpk} = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:526:5
			assign conv_target_q = 1'sb0;
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:529:3
	generate
		if ((DivSqrtSel != 2'd1) && !ExtRegEna) begin : genblk7
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:531:5
			assign simd_synch_rdy = (EnableVectors ? &divsqrt_ready[NUM_DIVSQRT_LANES - 1:0] : divsqrt_ready[0]);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:532:5
			assign simd_synch_done = (EnableVectors ? &divsqrt_done[NUM_DIVSQRT_LANES - 1:0] : divsqrt_done[0]);
		end
		else begin : genblk7
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:535:5
			assign simd_synch_rdy = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:536:5
			assign simd_synch_done = 1'sb0;
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:542:3
	assign {result_fmt_is_int, result_is_vector, result_fmt} = lane_aux[0+:AUX_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:544:3
	assign result_o = (result_fmt_is_int ? ifmt_slice_result[result_fmt * Width+:Width] : fmt_slice_result[result_fmt * Width+:Width]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:548:3
	assign extension_bit_o = lane_ext_bit[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:549:3
	assign tag_o = lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + 0+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:550:3
	assign busy_o = |lane_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:552:3
	assign out_valid_o = lane_out_valid[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:555:3
	always @(*) begin : output_processing
		// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:557:5
		reg [4:0] temp_status;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:558:5
		temp_status = 1'sb0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:559:5
		begin : sv2v_autoblock_12
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:559:10
			reg signed [31:0] i;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:559:10
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:560:7
					temp_status = temp_status | (lane_status[i * 5+:5] & {5 {lane_masks[i]}});
				end
		end
		// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_multifmt_slice.sv:561:5
		status_o = temp_status;
	end
endmodule
module fpnew_divsqrt_multi_68C3A_AC02A (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	dst_fmt_i,
	tag_i,
	mask_i,
	aux_i,
	vectorial_op_i,
	in_valid_i,
	in_ready_o,
	divsqrt_done_o,
	simd_synch_done_i,
	divsqrt_ready_o,
	simd_synch_rdy_i,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	mask_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o,
	reg_ena_i
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// removed localparam type TagType_TagType_TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:19:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:21:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:22:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:23:38
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:24:38
	// removed localparam type AuxType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:26:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:307:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:319:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:320:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:5
			begin : sv2v_autoblock_1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:323:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:27:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:28:14
	localparam [31:0] ExtRegEnaWidth = (NumPipeRegs == 0 ? 1 : NumPipeRegs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:30:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:31:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:33:3
	input wire [(2 * WIDTH) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:34:3
	input wire [9:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:35:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:36:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:37:3
	input wire [2:0] dst_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:38:3
	input wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:39:3
	input wire mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:40:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:41:3
	input wire vectorial_op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:43:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:44:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:45:3
	output wire divsqrt_done_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:46:3
	input wire simd_synch_done_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:47:3
	output wire divsqrt_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:48:3
	input wire simd_synch_rdy_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:49:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:51:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:52:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:53:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:54:3
	output wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:55:3
	output wire mask_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:56:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:58:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:59:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:61:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:63:3
	input wire [ExtRegEnaWidth - 1:0] reg_ena_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:70:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:75:3
	localparam NUM_OUT_REGS = ((PipeConfig == 2'd1) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:85:3
	wire [(2 * WIDTH) - 1:0] operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:86:3
	wire [2:0] rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:87:3
	wire [3:0] op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:88:3
	wire [2:0] dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:89:3
	wire in_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:92:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:93:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:94:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:95:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:96:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] inp_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:97:3
	reg [0:NUM_INP_REGS] inp_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:98:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:99:3
	reg [0:NUM_INP_REGS] inp_pipe_vec_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:100:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:102:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:105:3
	wire [2 * WIDTH:1] sv2v_tmp_83757;
	assign sv2v_tmp_83757 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_83757;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:106:3
	wire [3:1] sv2v_tmp_857E9;
	assign sv2v_tmp_857E9 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_857E9;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:107:3
	wire [4:1] sv2v_tmp_4BFFB;
	assign sv2v_tmp_4BFFB = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_4BFFB;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:108:3
	wire [3:1] sv2v_tmp_54055;
	assign sv2v_tmp_54055 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_54055;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:109:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_A168A;
	assign sv2v_tmp_A168A = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_A168A;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:110:3
	wire [1:1] sv2v_tmp_407DF;
	assign sv2v_tmp_407DF = mask_i;
	always @(*) inp_pipe_mask_q[0] = sv2v_tmp_407DF;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:111:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_51D85;
	assign sv2v_tmp_51D85 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_51D85;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:112:3
	wire [1:1] sv2v_tmp_EFF0C;
	assign sv2v_tmp_EFF0C = vectorial_op_i;
	always @(*) inp_pipe_vec_op_q[0] = sv2v_tmp_EFF0C;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:113:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:115:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:117:3
	genvar _gv_i_219;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] sv2v_cast_48BE4;
		input reg [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] inp;
		sv2v_cast_48BE4 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (_gv_i_219 = 0; _gv_i_219 < NUM_INP_REGS; _gv_i_219 = _gv_i_219 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_219;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:119:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:123:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:125:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:125:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:125:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:125:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:127:5
			assign reg_ena = (inp_pipe_ready[i] & inp_pipe_valid_q[i]) | reg_ena_i[i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:129:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:129:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:129:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:129:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:130:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:130:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:130:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:130:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:131:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:131:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:131:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:131:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:132:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:132:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:132:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:132:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:133:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:133:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:133:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:133:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:134:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:134:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:134:183
					inp_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:134:291
					inp_pipe_mask_q[i + 1] <= (reg_ena ? inp_pipe_mask_q[i] : inp_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:135:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:135:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:135:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:135:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:136:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:136:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:136:193
					inp_pipe_vec_op_q[i + 1] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:136:301
					inp_pipe_vec_op_q[i + 1] <= (reg_ena ? inp_pipe_vec_op_q[i] : inp_pipe_vec_op_q[i + 1]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:139:3
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:140:3
	assign rnd_mode_q = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:141:3
	assign op_q = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:142:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:143:3
	assign in_valid_q = inp_pipe_valid_q[NUM_INP_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:145:3
	reg ext_op_start_q;
	// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:146:55
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:146:111
		if (!rst_ni)
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:146:167
			ext_op_start_q <= 1'b0;
		else
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:146:275
			ext_op_start_q <= reg_ena_i[NUM_INP_REGS - 1];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:151:3
	reg [1:0] divsqrt_fmt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:152:3
	reg [127:0] divsqrt_operands;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:153:3
	reg input_is_fp8;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:156:3
	always @(*) begin : translate_fmt
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:157:5
		case (dst_fmt_q)
			sv2v_cast_0BC43('d0):
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:158:27
				divsqrt_fmt = 2'b00;
			sv2v_cast_0BC43('d1):
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:159:27
				divsqrt_fmt = 2'b01;
			sv2v_cast_0BC43('d2):
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:160:27
				divsqrt_fmt = 2'b10;
			sv2v_cast_0BC43('d4):
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:161:27
				divsqrt_fmt = 2'b11;
			default:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:162:27
				divsqrt_fmt = 2'b10;
		endcase
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:166:5
		input_is_fp8 = FpFmtConfig[sv2v_cast_0BC43('d3)] & (dst_fmt_q == sv2v_cast_0BC43('d3));
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:169:5
		divsqrt_operands[0+:64] = (input_is_fp8 ? operands_q[0+:WIDTH] << 8 : operands_q[0+:WIDTH]);
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:170:5
		divsqrt_operands[64+:64] = (input_is_fp8 ? operands_q[WIDTH+:WIDTH] << 8 : operands_q[WIDTH+:WIDTH]);
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:177:3
	reg in_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:178:3
	wire div_valid;
	wire sqrt_valid;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:179:3
	wire unit_ready;
	wire unit_done;
	reg unit_done_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:180:3
	wire op_starting;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:181:3
	reg out_valid;
	wire out_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:182:3
	reg unit_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:183:3
	wire simd_synch_done;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:185:3
	// removed localparam type fsm_state_e
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:186:3
	reg [1:0] state_q;
	reg [1:0] state_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:189:3
	assign div_valid = (((in_valid_q & in_ready) & ~flush_i) | ext_op_start_q) & (op_q == sv2v_cast_A53F3(4));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:190:3
	assign sqrt_valid = (((in_valid_q & in_ready) & ~flush_i) | ext_op_start_q) & (op_q != sv2v_cast_A53F3(4));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:191:3
	assign op_starting = div_valid | sqrt_valid;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:194:3
	reg result_is_fp8_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:195:3
	reg [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] result_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:196:3
	reg result_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:197:3
	reg [AuxType_AUX_BITS - 1:0] result_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:198:3
	reg result_vec_op_q;
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:201:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:201:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:201:182
			result_is_fp8_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:201:290
			result_is_fp8_q <= (op_starting ? input_is_fp8 : result_is_fp8_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:202:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:202:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:202:182
			result_tag_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:202:290
			result_tag_q <= (op_starting ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : result_tag_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:203:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:203:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:203:182
			result_mask_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:203:290
			result_mask_q <= (op_starting ? inp_pipe_mask_q[NUM_INP_REGS] : result_mask_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:204:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:204:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:204:182
			result_aux_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:204:290
			result_aux_q <= (op_starting ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : result_aux_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:205:73
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:205:129
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:205:185
			result_vec_op_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:205:293
			result_vec_op_q <= (op_starting ? inp_pipe_vec_op_q[NUM_INP_REGS] : result_vec_op_q);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:208:3
	assign simd_synch_done = simd_synch_done_i || ~result_vec_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:213:3
	wire unit_done_clear;
	// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:214:230
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:214:308
		if (!rst_ni)
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:214:386
			unit_done_q <= 1'b0;
		else
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:214:538
			unit_done_q <= (unit_done_clear ? 1'b0 : (unit_done ? unit_done : unit_done_q));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:215:3
	assign unit_done_clear = simd_synch_done | reg_ena_i[NUM_INP_REGS - 1];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:217:3
	assign divsqrt_done_o = (unit_done_q | unit_done) & result_vec_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:221:3
	assign divsqrt_ready_o = in_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:223:3
	assign inp_pipe_ready[NUM_INP_REGS] = (result_vec_op_q ? simd_synch_rdy_i : in_ready);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:226:3
	always @(*) begin : flag_fsm
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:228:5
		in_ready = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:229:5
		out_valid = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:230:5
		unit_busy = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:231:5
		state_d = state_q;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:233:5
		case (state_q)
			2'd0: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:236:9
				in_ready = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:237:9
				if (in_valid_q && unit_ready)
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:238:11
					state_d = 2'd1;
			end
			2'd1: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:243:9
				unit_busy = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:245:9
				if (simd_synch_done_i || (~result_vec_op_q && unit_done)) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:246:11
					out_valid = 1'b1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:248:11
					if (out_ready) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:249:13
						state_d = 2'd0;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:250:13
						in_ready = 1'b1;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:251:13
						if (in_valid_q && unit_ready)
							// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:252:15
							state_d = 2'd1;
					end
					else
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:256:13
						state_d = 2'd2;
				end
			end
			2'd2: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:262:9
				unit_busy = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:263:9
				out_valid = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:265:9
				if (out_ready) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:266:11
					state_d = 2'd0;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:267:11
					if (in_valid_q && unit_ready) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:268:13
						in_ready = 1'b1;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:269:13
						state_d = 2'd1;
					end
				end
			end
			default:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:274:16
				state_d = 2'd0;
		endcase
		if (flush_i) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:279:7
			unit_busy = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:280:7
			out_valid = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:281:7
			state_d = 2'd0;
		end
	end
	// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:286:30
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:286:86
		if (!rst_ni)
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:286:142
			state_q <= 2'd0;
		else
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:286:250
			state_q <= state_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:291:3
	wire [63:0] unit_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:292:3
	wire [WIDTH - 1:0] adjusted_result;
	reg [WIDTH - 1:0] held_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:293:3
	wire [4:0] unit_status;
	reg [4:0] held_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:294:3
	wire hold_en;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:296:3
	// removed localparam type sv2v_uu_i_divsqrt_lei_Precision_ctl_SI
	localparam [5:0] sv2v_uu_i_divsqrt_lei_ext_Precision_ctl_SI_0 = 1'sb0;
	div_sqrt_top_mvp i_divsqrt_lei(
		.Clk_CI(clk_i),
		.Rst_RBI(rst_ni),
		.Div_start_SI(div_valid),
		.Sqrt_start_SI(sqrt_valid),
		.Operand_a_DI(divsqrt_operands[0+:64]),
		.Operand_b_DI(divsqrt_operands[64+:64]),
		.RM_SI(rnd_mode_q),
		.Precision_ctl_SI(sv2v_uu_i_divsqrt_lei_ext_Precision_ctl_SI_0),
		.Format_sel_SI(divsqrt_fmt),
		.Kill_SI(flush_i | reg_ena_i[NUM_INP_REGS - 1]),
		.Result_DO(unit_result),
		.Fflags_SO(unit_status),
		.Ready_SO(unit_ready),
		.Done_SO(unit_done)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:314:3
	assign adjusted_result = (result_is_fp8_q ? unit_result >> 8 : unit_result);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:318:3
	assign hold_en = (unit_done & (~simd_synch_done_i | ~out_ready)) & ~(~result_vec_op_q & out_ready);
	// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:320:54
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:320:96
		held_result_q <= (hold_en ? adjusted_result : held_result_q);
	// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:321:54
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:321:96
		held_status_q <= (hold_en ? unit_status : held_status_q);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:326:3
	wire [WIDTH - 1:0] result_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:327:3
	wire [4:0] status_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:329:3
	assign result_d = (unit_done_q ? held_result_q : adjusted_result);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:330:3
	assign status_d = (unit_done_q ? held_status_q : unit_status);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:336:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:337:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:338:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] out_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:339:3
	reg [0:NUM_OUT_REGS] out_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:340:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:341:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:343:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:346:3
	wire [WIDTH * 1:1] sv2v_tmp_6C30D;
	assign sv2v_tmp_6C30D = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_6C30D;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:347:3
	wire [5:1] sv2v_tmp_2ED07;
	assign sv2v_tmp_2ED07 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_2ED07;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:348:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_D8454;
	assign sv2v_tmp_D8454 = result_tag_q;
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_D8454;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:349:3
	wire [1:1] sv2v_tmp_11413;
	assign sv2v_tmp_11413 = result_mask_q;
	always @(*) out_pipe_mask_q[0] = sv2v_tmp_11413;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:350:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_A8613;
	assign sv2v_tmp_A8613 = result_aux_q;
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_A8613;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:351:3
	wire [1:1] sv2v_tmp_D06FD;
	assign sv2v_tmp_D06FD = out_valid;
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_D06FD;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:353:3
	assign out_ready = out_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:355:3
	genvar _gv_i_220;
	generate
		for (_gv_i_220 = 0; _gv_i_220 < NUM_OUT_REGS; _gv_i_220 = _gv_i_220 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_220;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:357:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:361:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:363:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:363:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:363:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:363:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:365:5
			assign reg_ena = (out_pipe_ready[i] & out_pipe_valid_q[i]) | reg_ena_i[NUM_INP_REGS + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:367:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:367:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:367:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:367:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:368:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:368:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:368:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:368:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:369:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:369:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:369:189
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:369:297
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:370:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:370:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:370:179
					out_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:370:287
					out_pipe_mask_q[i + 1] <= (reg_ena ? out_pipe_mask_q[i] : out_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:371:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:371:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:371:189
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:371:297
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:374:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:376:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:377:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:378:3
	assign extension_bit_o = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:379:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:380:3
	assign mask_o = out_pipe_mask_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:381:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:382:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_multi.sv:383:3
	assign busy_o = |{inp_pipe_valid_q, unit_busy, out_pipe_valid_q};
endmodule
module fpnew_divsqrt_th_32_2BDD9_C9EC9 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	tag_i,
	mask_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	mask_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o,
	reg_ena_i
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// removed localparam type TagType_TagType_TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:24:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:25:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:26:38
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:27:38
	// removed localparam type AuxType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:29:14
	localparam [31:0] WIDTH = 32;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:30:14
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:31:14
	localparam [31:0] ExtRegEnaWidth = (NumPipeRegs == 0 ? 1 : NumPipeRegs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:33:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:34:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:36:3
	input wire [63:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:37:3
	input wire [9:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:38:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:39:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:40:3
	input wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:41:3
	input wire mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:42:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:44:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:45:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:46:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:48:3
	output wire [31:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:49:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:50:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:51:3
	output wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:52:3
	output wire mask_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:53:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:55:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:56:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:58:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:60:3
	input wire [ExtRegEnaWidth - 1:0] reg_ena_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:67:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:72:3
	localparam NUM_OUT_REGS = ((PipeConfig == 2'd1) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:82:3
	wire [63:0] operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:83:3
	wire [2:0] rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:84:3
	wire [3:0] op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:85:3
	wire in_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:88:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * 32) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * 32) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * 32) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * 32) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * 32 : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * 32)] inp_pipe_operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:89:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:90:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:91:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] inp_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:92:3
	reg [0:NUM_INP_REGS] inp_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:93:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:94:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:96:3
	reg [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:99:3
	wire [64:1] sv2v_tmp_6F41F;
	assign sv2v_tmp_6F41F = operands_i;
	always @(*) inp_pipe_operands_q[32 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:64] = sv2v_tmp_6F41F;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:100:3
	wire [3:1] sv2v_tmp_CE431;
	assign sv2v_tmp_CE431 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_CE431;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:101:3
	wire [4:1] sv2v_tmp_B00A7;
	assign sv2v_tmp_B00A7 = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_B00A7;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:102:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_B7AFE;
	assign sv2v_tmp_B7AFE = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_B7AFE;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:103:3
	wire [1:1] sv2v_tmp_407DF;
	assign sv2v_tmp_407DF = mask_i;
	always @(*) inp_pipe_mask_q[0] = sv2v_tmp_407DF;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:104:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_49B77;
	assign sv2v_tmp_49B77 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_49B77;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:105:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:107:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:109:3
	genvar _gv_i_221;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] sv2v_cast_48BE4;
		input reg [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] inp;
		sv2v_cast_48BE4 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (_gv_i_221 = 0; _gv_i_221 < NUM_INP_REGS; _gv_i_221 = _gv_i_221 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_221;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:111:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:115:5
			wire [1:1] sv2v_tmp_2ABCB;
			assign sv2v_tmp_2ABCB = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			always @(*) inp_pipe_ready[i] = sv2v_tmp_2ABCB;
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:117:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:117:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:117:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:117:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:119:5
			assign reg_ena = (inp_pipe_ready[i] & inp_pipe_valid_q[i]) | reg_ena_i[i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:121:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:121:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:121:183
					inp_pipe_operands_q[32 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:64] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:121:291
					inp_pipe_operands_q[32 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:64] <= (reg_ena ? inp_pipe_operands_q[32 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:64] : inp_pipe_operands_q[32 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:64]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:122:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:122:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:122:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:122:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:123:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:123:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:123:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:123:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:124:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:124:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:124:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:124:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:125:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:125:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:125:183
					inp_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:125:291
					inp_pipe_mask_q[i + 1] <= (reg_ena ? inp_pipe_mask_q[i] : inp_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:126:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:126:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:126:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:126:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:129:3
	assign operands_q = inp_pipe_operands_q[32 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:64];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:130:3
	assign rnd_mode_q = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:131:3
	assign op_q = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:132:3
	assign in_valid_q = inp_pipe_valid_q[NUM_INP_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:137:3
	reg in_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:138:3
	wire div_op;
	wire sqrt_op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:139:3
	reg unit_ready_q;
	reg unit_done;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:140:3
	wire op_starting;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:141:3
	reg out_valid;
	wire out_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:142:3
	reg hold_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:143:3
	reg data_is_held;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:144:3
	reg unit_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:146:3
	// removed localparam type fsm_state_e
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:147:3
	reg [1:0] state_q;
	reg [1:0] state_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:150:3
	assign div_op = ((in_valid_q & (op_q == sv2v_cast_A53F3(4))) & in_ready) & ~flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:151:3
	assign sqrt_op = ((in_valid_q & (op_q == sv2v_cast_A53F3(5))) & in_ready) & ~flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:152:3
	assign op_starting = div_op | sqrt_op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:154:3
	wire fdsu_fpu_ex1_stall;
	reg fdsu_fpu_ex1_stall_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:155:3
	wire div_op_d;
	reg div_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:156:3
	wire sqrt_op_d;
	reg sqrt_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:158:3
	assign div_op_d = (fdsu_fpu_ex1_stall ? div_op : 1'b0);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:159:3
	assign sqrt_op_d = (fdsu_fpu_ex1_stall ? sqrt_op : 1'b0);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:161:58
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:161:114
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:161:170
			fdsu_fpu_ex1_stall_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:161:278
			fdsu_fpu_ex1_stall_q <= fdsu_fpu_ex1_stall;
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:162:36
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:162:92
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:162:148
			div_op_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:162:256
			div_op_q <= div_op_d;
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:163:38
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:163:94
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:163:150
			sqrt_op_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:163:258
			sqrt_op_q <= sqrt_op_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:166:3
	always @(*) begin : flag_fsm
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:168:5
		in_ready = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:169:5
		out_valid = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:170:5
		hold_result = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:171:5
		data_is_held = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:172:5
		unit_busy = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:173:5
		state_d = state_q;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:174:5
		inp_pipe_ready[NUM_INP_REGS] = unit_ready_q;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:176:5
		case (state_q)
			2'd0: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:180:9
				in_ready = unit_ready_q;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:181:9
				if (in_valid_q && unit_ready_q) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:182:11
					inp_pipe_ready[NUM_INP_REGS] = unit_ready_q && !fdsu_fpu_ex1_stall;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:183:11
					state_d = 2'd1;
				end
			end
			2'd1: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:188:9
				inp_pipe_ready[NUM_INP_REGS] = fdsu_fpu_ex1_stall_q;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:189:9
				unit_busy = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:191:9
				if (unit_done) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:192:11
					out_valid = 1'b1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:194:11
					if (out_ready) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:195:13
						state_d = 2'd0;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:196:13
						if (in_valid_q && unit_ready_q) begin
							// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:197:15
							in_ready = 1'b1;
							// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:198:15
							state_d = 2'd1;
						end
					end
					else begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:202:13
						hold_result = 1'b1;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:203:13
						state_d = 2'd2;
					end
				end
			end
			2'd2: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:209:9
				unit_busy = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:210:9
				data_is_held = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:211:9
				out_valid = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:213:9
				if (out_ready) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:214:11
					state_d = 2'd0;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:215:11
					if (in_valid_q && unit_ready_q) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:216:13
						in_ready = 1'b1;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:217:13
						state_d = 2'd1;
					end
				end
			end
			default:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:222:16
				state_d = 2'd0;
		endcase
		if (flush_i) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:227:7
			unit_busy = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:228:7
			out_valid = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:229:7
			state_d = 2'd0;
		end
	end
	// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:234:30
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:234:86
		if (!rst_ni)
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:234:142
			state_q <= 2'd0;
		else
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:234:250
			state_q <= state_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:237:3
	reg [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] result_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:238:3
	reg [AuxType_AUX_BITS - 1:0] result_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:239:3
	reg result_mask_q;
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:242:69
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:242:125
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:242:181
			result_tag_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:242:289
			result_tag_q <= (op_starting ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : result_tag_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:243:69
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:243:125
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:243:181
			result_mask_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:243:289
			result_mask_q <= (op_starting ? inp_pipe_mask_q[NUM_INP_REGS] : result_mask_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:244:69
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:244:125
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:244:181
			result_aux_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:244:289
			result_aux_q <= (op_starting ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : result_aux_q);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:249:3
	reg [31:0] unit_result;
	reg [31:0] held_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:250:3
	reg [4:0] unit_status;
	reg [4:0] held_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:253:3
	reg ctrl_fdsu_ex1_sel;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:254:3
	wire fdsu_fpu_ex1_cmplt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:255:3
	wire [4:0] fdsu_fpu_ex1_fflags;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:256:3
	wire [7:0] fdsu_fpu_ex1_special_sel;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:257:3
	wire [3:0] fdsu_fpu_ex1_special_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:258:3
	wire fdsu_fpu_no_op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:259:3
	reg [2:0] idu_fpu_ex1_eu_sel;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:260:3
	wire [31:0] fdsu_frbus_data;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:261:3
	wire [4:0] fdsu_frbus_fflags;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:262:3
	wire fdsu_frbus_wb_vld;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:265:3
	wire [31:0] dp_frbus_ex2_data;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:266:3
	wire [4:0] dp_frbus_ex2_fflags;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:267:3
	wire [2:0] dp_xx_ex1_cnan;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:268:3
	wire [2:0] dp_xx_ex1_id;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:269:3
	wire [2:0] dp_xx_ex1_inf;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:270:3
	wire [2:0] dp_xx_ex1_norm;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:271:3
	wire [2:0] dp_xx_ex1_qnan;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:272:3
	wire [2:0] dp_xx_ex1_snan;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:273:3
	wire [2:0] dp_xx_ex1_zero;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:274:3
	wire ex2_inst_wb;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:275:3
	wire ex2_inst_wb_vld_d;
	reg ex2_inst_wb_vld_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:278:3
	wire [31:0] fpu_idu_fwd_data;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:279:3
	wire [4:0] fpu_idu_fwd_fflags;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:280:3
	wire fpu_idu_fwd_vld;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:282:3
	reg unit_ready_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:285:3
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:286:5
		if (op_starting && unit_ready_q) begin
			begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:287:7
				if (ex2_inst_wb && ex2_inst_wb_vld_q)
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:288:9
					unit_ready_d = 1'b1;
				else
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:290:9
					unit_ready_d = 1'b0;
			end
		end
		else if (fpu_idu_fwd_vld | flush_i)
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:293:7
			unit_ready_d = 1'b1;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:295:7
			unit_ready_d = unit_ready_q;
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:299:46
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:299:102
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:299:158
			unit_ready_q <= 1'b1;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:299:266
			unit_ready_q <= unit_ready_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:302:3
	always @(*) begin
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:303:5
		ctrl_fdsu_ex1_sel = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:304:5
		idu_fpu_ex1_eu_sel = 3'h0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:305:5
		if (op_starting) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:306:7
			ctrl_fdsu_ex1_sel = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:307:7
			idu_fpu_ex1_eu_sel = 3'h4;
		end
		else if (fdsu_fpu_ex1_stall_q) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:309:7
			ctrl_fdsu_ex1_sel = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:310:7
			idu_fpu_ex1_eu_sel = 3'h4;
		end
		else begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:312:7
			ctrl_fdsu_ex1_sel = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:313:7
			idu_fpu_ex1_eu_sel = 3'h0;
		end
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:317:3
	pa_fdsu_top i_divsqrt_thead(
		.cp0_fpu_icg_en(1'b0),
		.cp0_fpu_xx_dqnan(1'b0),
		.cp0_yy_clk_en(1'b1),
		.cpurst_b(rst_ni),
		.ctrl_fdsu_ex1_sel(ctrl_fdsu_ex1_sel),
		.ctrl_xx_ex1_cmplt_dp(ctrl_fdsu_ex1_sel),
		.ctrl_xx_ex1_inst_vld(ctrl_fdsu_ex1_sel),
		.ctrl_xx_ex1_stall(fdsu_fpu_ex1_stall),
		.ctrl_xx_ex1_warm_up(1'b0),
		.ctrl_xx_ex2_warm_up(1'b0),
		.ctrl_xx_ex3_warm_up(1'b0),
		.dp_xx_ex1_cnan(dp_xx_ex1_cnan),
		.dp_xx_ex1_id(dp_xx_ex1_id),
		.dp_xx_ex1_inf(dp_xx_ex1_inf),
		.dp_xx_ex1_qnan(dp_xx_ex1_qnan),
		.dp_xx_ex1_rm(rnd_mode_q),
		.dp_xx_ex1_snan(dp_xx_ex1_snan),
		.dp_xx_ex1_zero(dp_xx_ex1_zero),
		.fdsu_fpu_debug_info(),
		.fdsu_fpu_ex1_cmplt(fdsu_fpu_ex1_cmplt),
		.fdsu_fpu_ex1_cmplt_dp(),
		.fdsu_fpu_ex1_fflags(fdsu_fpu_ex1_fflags),
		.fdsu_fpu_ex1_special_sel(fdsu_fpu_ex1_special_sel),
		.fdsu_fpu_ex1_special_sign(fdsu_fpu_ex1_special_sign),
		.fdsu_fpu_ex1_stall(fdsu_fpu_ex1_stall),
		.fdsu_fpu_no_op(fdsu_fpu_no_op),
		.fdsu_frbus_data(fdsu_frbus_data),
		.fdsu_frbus_fflags(fdsu_frbus_fflags),
		.fdsu_frbus_freg(),
		.fdsu_frbus_wb_vld(fdsu_frbus_wb_vld),
		.forever_cpuclk(clk_i),
		.frbus_fdsu_wb_grant(fdsu_frbus_wb_vld),
		.idu_fpu_ex1_dst_freg(5'h0f),
		.idu_fpu_ex1_eu_sel(idu_fpu_ex1_eu_sel),
		.idu_fpu_ex1_func({8'b00000000, div_op | div_op_q, sqrt_op | sqrt_op_q}),
		.idu_fpu_ex1_srcf0(operands_q[31-:32]),
		.idu_fpu_ex1_srcf1(operands_q[63-:32]),
		.pad_yy_icg_scan_en(1'b0),
		.rtu_xx_ex1_cancel(1'b0),
		.rtu_xx_ex2_cancel(1'b0),
		.rtu_yy_xx_async_flush(flush_i),
		.rtu_yy_xx_flush(1'b0)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:362:3
	pa_fpu_dp x_pa_fpu_dp(
		.cp0_fpu_icg_en(1'b0),
		.cp0_fpu_xx_rm(rnd_mode_q),
		.cp0_yy_clk_en(1'b1),
		.ctrl_xx_ex1_inst_vld(ctrl_fdsu_ex1_sel),
		.ctrl_xx_ex1_stall(1'b0),
		.ctrl_xx_ex1_warm_up(1'b0),
		.dp_frbus_ex2_data(dp_frbus_ex2_data),
		.dp_frbus_ex2_fflags(dp_frbus_ex2_fflags),
		.dp_xx_ex1_cnan(dp_xx_ex1_cnan),
		.dp_xx_ex1_id(dp_xx_ex1_id),
		.dp_xx_ex1_inf(dp_xx_ex1_inf),
		.dp_xx_ex1_norm(dp_xx_ex1_norm),
		.dp_xx_ex1_qnan(dp_xx_ex1_qnan),
		.dp_xx_ex1_snan(dp_xx_ex1_snan),
		.dp_xx_ex1_zero(dp_xx_ex1_zero),
		.ex2_inst_wb(ex2_inst_wb),
		.fdsu_fpu_ex1_fflags(fdsu_fpu_ex1_fflags),
		.fdsu_fpu_ex1_special_sel(fdsu_fpu_ex1_special_sel),
		.fdsu_fpu_ex1_special_sign(fdsu_fpu_ex1_special_sign),
		.forever_cpuclk(clk_i),
		.idu_fpu_ex1_eu_sel(idu_fpu_ex1_eu_sel),
		.idu_fpu_ex1_func({8'b00000000, div_op, sqrt_op}),
		.idu_fpu_ex1_gateclk_vld(fdsu_fpu_ex1_cmplt),
		.idu_fpu_ex1_rm(rnd_mode_q),
		.idu_fpu_ex1_srcf0(operands_q[31-:32]),
		.idu_fpu_ex1_srcf1(operands_q[63-:32]),
		.idu_fpu_ex1_srcf2(1'sb0),
		.pad_yy_icg_scan_en(1'b0)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:393:3
	assign ex2_inst_wb_vld_d = ctrl_fdsu_ex1_sel;
	// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:394:48
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:394:104
		if (!rst_ni)
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:394:160
			ex2_inst_wb_vld_q <= 1'sb0;
		else
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:394:268
			ex2_inst_wb_vld_q <= ex2_inst_wb_vld_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:396:3
	pa_fpu_frbus x_pa_fpu_frbus(
		.ctrl_frbus_ex2_wb_req(ex2_inst_wb & ex2_inst_wb_vld_q),
		.dp_frbus_ex2_data(dp_frbus_ex2_data),
		.dp_frbus_ex2_fflags(dp_frbus_ex2_fflags),
		.fdsu_frbus_data(fdsu_frbus_data),
		.fdsu_frbus_fflags(fdsu_frbus_fflags),
		.fdsu_frbus_wb_vld(fdsu_frbus_wb_vld),
		.fpu_idu_fwd_data(fpu_idu_fwd_data),
		.fpu_idu_fwd_fflags(fpu_idu_fwd_fflags),
		.fpu_idu_fwd_vld(fpu_idu_fwd_vld)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:408:3
	always @(*) begin
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:409:5
		unit_result[31:0] = fpu_idu_fwd_data[31:0];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:410:5
		unit_status[4:0] = fpu_idu_fwd_fflags[4:0];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:411:5
		unit_done = fpu_idu_fwd_vld;
	end
	// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:415:54
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:415:96
		held_result_q <= (hold_result ? unit_result : held_result_q);
	// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:416:54
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:416:96
		held_status_q <= (hold_result ? unit_status : held_status_q);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:421:3
	wire [31:0] result_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:422:3
	wire [4:0] status_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:424:3
	assign result_d = (data_is_held ? held_result_q : unit_result);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:425:3
	assign status_d = (data_is_held ? held_status_q : unit_status);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:431:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:432:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:433:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] out_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:434:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:435:3
	reg [0:NUM_OUT_REGS] out_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:436:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:438:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:441:3
	wire [32:1] sv2v_tmp_37F39;
	assign sv2v_tmp_37F39 = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_37F39;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:442:3
	wire [5:1] sv2v_tmp_83427;
	assign sv2v_tmp_83427 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_83427;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:443:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_9961C;
	assign sv2v_tmp_9961C = result_tag_q;
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_9961C;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:444:3
	wire [1:1] sv2v_tmp_11413;
	assign sv2v_tmp_11413 = result_mask_q;
	always @(*) out_pipe_mask_q[0] = sv2v_tmp_11413;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:445:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_FA16D;
	assign sv2v_tmp_FA16D = result_aux_q;
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_FA16D;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:446:3
	wire [1:1] sv2v_tmp_D06FD;
	assign sv2v_tmp_D06FD = out_valid;
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_D06FD;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:448:3
	assign out_ready = out_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:450:3
	genvar _gv_i_222;
	generate
		for (_gv_i_222 = 0; _gv_i_222 < NUM_OUT_REGS; _gv_i_222 = _gv_i_222 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_222;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:452:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:456:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:458:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:458:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:458:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:458:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:460:5
			assign reg_ena = (out_pipe_ready[i] & out_pipe_valid_q[i]) | reg_ena_i[NUM_INP_REGS + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:462:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:462:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:462:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:462:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:463:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:463:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:463:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:463:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:464:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:464:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:464:189
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:464:297
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:465:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:465:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:465:179
					out_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:465:287
					out_pipe_mask_q[i + 1] <= (reg_ena ? out_pipe_mask_q[i] : out_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:466:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:466:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:466:189
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:466:297
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:469:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:471:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:472:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:473:3
	assign extension_bit_o = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:474:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:475:3
	assign mask_o = out_pipe_mask_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:476:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:477:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_32.sv:478:3
	assign busy_o = |{inp_pipe_valid_q, unit_busy, out_pipe_valid_q};
endmodule
module fpnew_fma_multi_6D055_6E71C (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	src2_fmt_i,
	dst_fmt_i,
	tag_i,
	mask_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	mask_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o,
	reg_ena_i
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// removed localparam type TagType_TagType_TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:19:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:20:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:21:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:22:38
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:23:38
	// removed localparam type AuxType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:25:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:307:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:319:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:320:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:5
			begin : sv2v_autoblock_1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:323:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:26:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:27:14
	localparam [31:0] ExtRegEnaWidth = (NumPipeRegs == 0 ? 1 : NumPipeRegs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:29:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:30:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:32:3
	input wire [(3 * WIDTH) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:33:3
	input wire [14:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:34:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:35:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:36:3
	input wire op_mod_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:37:3
	input wire [2:0] src_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:38:3
	input wire [2:0] src2_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:39:3
	input wire [2:0] dst_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:40:3
	input wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:41:3
	input wire mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:42:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:44:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:45:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:46:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:48:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:49:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:50:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:51:3
	output wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:52:3
	output wire mask_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:53:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:55:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:56:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:58:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:60:3
	input wire [ExtRegEnaWidth - 1:0] reg_ena_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:67:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:337:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:338:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:342:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:343:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:351:49
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:352:5
		reg [63:0] res;
		begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:353:5
			res = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:354:5
			begin : sv2v_autoblock_2
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:354:10
				reg [31:0] fmt;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:354:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:356:9
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt))));
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:357:9
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:69:3
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:70:3
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:73:3
	localparam [31:0] PRECISION_BITS = SUPER_MAN_BITS + 1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:75:3
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:76:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:80:3
	localparam [31:0] EXP_WIDTH = fpnew_pkg_maximum(SUPER_EXP_BITS + 2, LZC_RESULT_WIDTH);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:82:3
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 5);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:84:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:89:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:94:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:103:3
	// removed localparam type fp_t
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:113:3
	wire [(3 * WIDTH) - 1:0] operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:114:3
	wire [2:0] src_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:115:3
	wire [2:0] src2_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:116:3
	wire [2:0] dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:119:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:120:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)) + 1) * 3) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)) + 1) * 3) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3 : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3)] inp_pipe_is_boxed_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:121:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:122:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:123:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:124:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:125:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src2_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:126:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:127:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] inp_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:128:3
	reg [0:NUM_INP_REGS] inp_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:129:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:130:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:132:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:135:3
	wire [3 * WIDTH:1] sv2v_tmp_5DCC9;
	assign sv2v_tmp_5DCC9 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_5DCC9;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:136:3
	wire [15:1] sv2v_tmp_7F60B;
	assign sv2v_tmp_7F60B = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] = sv2v_tmp_7F60B;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:137:3
	wire [3:1] sv2v_tmp_700C1;
	assign sv2v_tmp_700C1 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_700C1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:138:3
	wire [4:1] sv2v_tmp_3923B;
	assign sv2v_tmp_3923B = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_3923B;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:139:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:140:3
	wire [3:1] sv2v_tmp_6B115;
	assign sv2v_tmp_6B115 = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_6B115;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:141:3
	wire [3:1] sv2v_tmp_539CB;
	assign sv2v_tmp_539CB = src2_fmt_i;
	always @(*) inp_pipe_src2_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_539CB;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:142:3
	wire [3:1] sv2v_tmp_B8677;
	assign sv2v_tmp_B8677 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_B8677;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:143:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_77526;
	assign sv2v_tmp_77526 = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_77526;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:144:3
	wire [1:1] sv2v_tmp_407DF;
	assign sv2v_tmp_407DF = mask_i;
	always @(*) inp_pipe_mask_q[0] = sv2v_tmp_407DF;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:145:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_129B7;
	assign sv2v_tmp_129B7 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_129B7;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:146:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:148:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:150:3
	genvar _gv_i_223;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] sv2v_cast_48BE4;
		input reg [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] inp;
		sv2v_cast_48BE4 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (_gv_i_223 = 0; _gv_i_223 < NUM_INP_REGS; _gv_i_223 = _gv_i_223 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_223;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:152:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:156:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:158:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:158:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:158:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:158:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:160:5
			assign reg_ena = (inp_pipe_ready[i] & inp_pipe_valid_q[i]) | reg_ena_i[i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:162:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:162:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:162:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:162:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:163:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:163:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:163:183
					inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:163:291
					inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= (reg_ena ? inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] : inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:164:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:164:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:164:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:164:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:165:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:165:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:165:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:165:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:166:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:166:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:166:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:166:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:167:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:167:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:167:207
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:167:315
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:168:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:168:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:168:207
					inp_pipe_src2_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:168:315
					inp_pipe_src2_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_src2_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_src2_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:169:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:169:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:169:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:169:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:170:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:170:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:170:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:170:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:171:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:171:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:171:183
					inp_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:171:291
					inp_pipe_mask_q[i + 1] <= (reg_ena ? inp_pipe_mask_q[i] : inp_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:172:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:172:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:172:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:172:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:175:3
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:176:3
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:177:3
	assign src2_fmt_q = inp_pipe_src2_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:178:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:183:3
	wire [14:0] fmt_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:184:3
	wire signed [(15 * SUPER_EXP_BITS) - 1:0] fmt_exponent;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:185:3
	wire [(15 * SUPER_MAN_BITS) - 1:0] fmt_mantissa;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:187:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [119:0] info_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:190:3
	genvar _gv_fmt_5;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic signed [SUPER_EXP_BITS - 1:0] sv2v_cast_A3BB6_signed;
		input reg signed [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_A3BB6_signed = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_52F63;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_52F63 = inp;
	endfunction
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_fmt_5 = 0; _gv_fmt_5 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_5 = _gv_fmt_5 + 1) begin : fmt_init_inputs
			localparam fmt = _gv_fmt_5;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:192:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:193:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:194:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:197:7
				localparam [2:0] FpFormat = sv2v_cast_0BC43(fmt);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:198:7
				wire [(3 * FP_WIDTH) - 1:0] trimmed_ops;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:201:7
				fpnew_classifier #(
					.FpFormat(FpFormat),
					.NumOperands(3)
				) i_fpnew_classifier(
					.operands_i(trimmed_ops),
					.is_boxed_i(inp_pipe_is_boxed_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1))) * 3+:3]),
					.info_o(info_q[8 * (fmt * 3)+:24])
				);
				genvar _gv_op_2;
				for (_gv_op_2 = 0; _gv_op_2 < 3; _gv_op_2 = _gv_op_2 + 1) begin : gen_operands
					localparam op = _gv_op_2;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:210:9
					assign trimmed_ops[op * fpnew_pkg_fp_width(sv2v_cast_0BC43(_gv_fmt_5))+:fpnew_pkg_fp_width(sv2v_cast_0BC43(_gv_fmt_5))] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH];
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:211:9
					assign fmt_sign[(fmt * 3) + op] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)];
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:212:9
					assign fmt_exponent[((fmt * 3) + op) * SUPER_EXP_BITS+:SUPER_EXP_BITS] = $signed({1'b0, operands_q[(op * WIDTH) + MAN_BITS+:EXP_BITS]});
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:213:9
					assign fmt_mantissa[((fmt * 3) + op) * SUPER_MAN_BITS+:SUPER_MAN_BITS] = {info_q[(((fmt * 3) + op) * 8) + 7], operands_q[(op * WIDTH) + (MAN_BITS - 1)-:MAN_BITS]} << (SUPER_MAN_BITS - MAN_BITS);
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:217:7
				assign info_q[8 * (fmt * 3)+:24] = {3 {sv2v_cast_8(fpnew_pkg_DONT_CARE)}};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:218:7
				assign fmt_sign[fmt * 3+:3] = fpnew_pkg_DONT_CARE;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:219:7
				assign fmt_exponent[SUPER_EXP_BITS * (fmt * 3)+:SUPER_EXP_BITS * 3] = {3 {sv2v_cast_A3BB6_signed(fpnew_pkg_DONT_CARE)}};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:220:7
				assign fmt_mantissa[SUPER_MAN_BITS * (fmt * 3)+:SUPER_MAN_BITS * 3] = {3 {sv2v_cast_52F63(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:224:3
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_a;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_b;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_c;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:225:3
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:239:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:347:40
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:348:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_A3BB6;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_A3BB6 = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_FC661;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_FC661 = inp;
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_705CC;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_705CC = inp;
	endfunction
	always @(*) begin : op_select
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:242:5
		operand_a = {fmt_sign[src_fmt_q * 3], fmt_exponent[(src_fmt_q * 3) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[(src_fmt_q * 3) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:243:5
		operand_b = {fmt_sign[(src_fmt_q * 3) + 1], fmt_exponent[((src_fmt_q * 3) + 1) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((src_fmt_q * 3) + 1) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:244:5
		operand_c = {fmt_sign[(src2_fmt_q * 3) + 2], fmt_exponent[((src2_fmt_q * 3) + 2) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((src2_fmt_q * 3) + 2) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:245:5
		info_a = info_q[(src_fmt_q * 3) * 8+:8];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:246:5
		info_b = info_q[((src_fmt_q * 3) + 1) * 8+:8];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:247:5
		info_c = info_q[((src2_fmt_q * 3) + 2) * 8+:8];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:250:5
		operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:252:5
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(0):
				;
			sv2v_cast_A53F3(1):
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:254:26
				operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = ~operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
			sv2v_cast_A53F3(2), sv2v_cast_A53F3(15): begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:257:9
				operand_a = {1'b0, sv2v_cast_A3BB6(fpnew_pkg_bias(src_fmt_q)), sv2v_cast_FC661(1'sb0)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:258:9
				info_a = 8'b10000001;
			end
			sv2v_cast_A53F3(3): begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:261:9
				if (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3] == 3'b010)
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:262:11
					operand_c = {1'b0, sv2v_cast_705CC(1'sb0), sv2v_cast_FC661(1'sb0)};
				else
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:264:11
					operand_c = {1'b1, sv2v_cast_705CC(1'sb0), sv2v_cast_FC661(1'sb0)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:265:9
				info_c = 8'b00100001;
			end
			default: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:268:9
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:269:9
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:270:9
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:271:9
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:272:9
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:273:9
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:281:3
	wire any_operand_inf;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:282:3
	wire any_operand_nan;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:283:3
	wire signalling_nan;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:284:3
	wire effective_subtraction;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:285:3
	wire tentative_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:288:3
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:289:3
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:290:3
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:292:3
	assign effective_subtraction = (operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))]) ^ operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:294:3
	assign tentative_sign = operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:299:3
	wire [WIDTH - 1:0] special_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:300:3
	wire [4:0] special_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:301:3
	wire result_is_special;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:303:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:304:3
	reg [24:0] fmt_special_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:305:3
	reg [4:0] fmt_result_is_special;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:308:3
	genvar _gv_fmt_6;
	generate
		for (_gv_fmt_6 = 0; _gv_fmt_6 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_6 = _gv_fmt_6 + 1) begin : gen_special_results
			localparam fmt = _gv_fmt_6;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:310:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:311:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:312:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:314:5
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:315:5
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:316:5
			localparam [MAN_BITS - 1:0] ZERO_MANTISSA = 1'sb0;
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:319:7
				always @(*) begin : special_results
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:320:9
					reg [FP_WIDTH - 1:0] special_res;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:323:9
					special_res = {1'b0, QNAN_EXPONENT, QNAN_MANTISSA};
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:324:9
					fmt_special_status[fmt * 5+:5] = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:325:9
					fmt_result_is_special[fmt] = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:331:9
					if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:332:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:333:11
						fmt_special_status[(fmt * 5) + 4] = 1'b1;
					end
					else if (any_operand_nan) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:336:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:337:11
						fmt_special_status[(fmt * 5) + 4] = signalling_nan;
					end
					else if (any_operand_inf) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:340:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:342:11
						if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
							// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:343:13
							fmt_special_status[(fmt * 5) + 4] = 1'b1;
						else if (info_a[4] || info_b[4])
							// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:347:13
							special_res = {operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
						else if (info_c[4])
							// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:351:13
							special_res = {operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
					end
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:355:9
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:356:9
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:359:7
				wire [WIDTH * 1:1] sv2v_tmp_7740B;
				assign sv2v_tmp_7740B = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_7740B;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:360:7
				wire [5:1] sv2v_tmp_899F4;
				assign sv2v_tmp_899F4 = 1'sb0;
				always @(*) fmt_special_status[fmt * 5+:5] = sv2v_tmp_899F4;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:361:7
				wire [1:1] sv2v_tmp_77BE5;
				assign sv2v_tmp_77BE5 = 1'b0;
				always @(*) fmt_result_is_special[fmt] = sv2v_tmp_77BE5;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:366:3
	assign result_is_special = fmt_result_is_special[dst_fmt_q];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:368:3
	assign special_status = fmt_special_status[dst_fmt_q * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:370:3
	assign special_result = fmt_special_result[dst_fmt_q * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:375:3
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:376:3
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:377:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:380:3
	assign exponent_a = $signed({1'b0, operand_a[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:381:3
	assign exponent_b = $signed({1'b0, operand_b[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:382:3
	assign exponent_c = $signed({1'b0, operand_c[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:386:3
	assign exponent_addend = (info_c[5] ? 1 : $signed(((exponent_c + $signed({1'b0, ~info_c[7]})) - $signed(fpnew_pkg_bias(src2_fmt_q))) + $signed(fpnew_pkg_bias(dst_fmt_q))));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:391:3
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(fpnew_pkg_bias(dst_fmt_q)) : $signed(((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - (2 * $signed(fpnew_pkg_bias(src_fmt_q)))) + $signed(fpnew_pkg_bias(dst_fmt_q))));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:398:3
	assign exponent_difference = exponent_addend - exponent_product;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:401:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:403:3
	always @(*) begin : addend_shift_amount
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:405:5
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:406:7
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:409:7
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:412:7
			addend_shamt = 0;
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:416:3
	wire [$clog2(SUPER_MAN_BITS) - 1:0] addend_lzc_count;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:417:3
	wire [$clog2(SUPER_MAN_BITS):0] addend_lzc_count_sgn;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:418:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_normalize_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:421:3
	lzc #(
		.WIDTH(SUPER_MAN_BITS),
		.MODE(1)
	) i_addend_lzc(
		.in_i(operand_c[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]),
		.cnt_o(addend_lzc_count),
		.empty_o()
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:430:3
	assign addend_lzc_count_sgn = $signed({1'b0, addend_lzc_count});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:433:3
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:435:5
		if (info_c[7] || info_c[5])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:436:7
			addend_normalize_shamt = 0;
		else if (exponent_addend <= 1)
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:439:7
			addend_normalize_shamt = 0;
		else if ((addend_lzc_count_sgn + 1) < exponent_addend)
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:442:7
			addend_normalize_shamt = addend_lzc_count + 1;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:445:7
			addend_normalize_shamt = exponent_addend - 1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:450:3
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend - addend_normalize_shamt : exponent_product);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:455:3
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:456:3
	wire [(2 * PRECISION_BITS) - 1:0] product;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:457:3
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:460:3
	assign mantissa_a = {info_a[7], operand_a[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:461:3
	assign mantissa_b = {info_b[7], operand_b[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:462:3
	assign mantissa_c = {info_c[7], operand_c[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:465:3
	assign product = mantissa_a * mantissa_b;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:470:3
	assign product_shifted = product << 2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:475:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:476:3
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:477:3
	wire sticky_before_add;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:478:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:479:3
	wire inject_carry_in;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:489:3
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:492:3
	assign sticky_before_add = |addend_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:495:3
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:496:3
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:501:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_pos;
	wire [(3 * PRECISION_BITS) + 4:0] sum_neg;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:502:3
	wire sum_carry;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:503:3
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:504:3
	wire final_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:507:3
	assign sum_pos = (product_shifted + addend_shifted) + inject_carry_in;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:508:3
	assign sum_carry = sum_pos[(3 * PRECISION_BITS) + 4];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:513:3
	assign sum_neg = addend_after_shift - product_shifted;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:516:3
	assign sum = (effective_subtraction && ~sum_carry ? sum_neg : sum_pos);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:519:3
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:527:3
	wire effective_subtraction_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:528:3
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:529:3
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:530:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:531:3
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:532:3
	wire sticky_before_add_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:533:3
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:534:3
	wire final_sign_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:535:3
	wire [2:0] dst_fmt_q2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:536:3
	wire [2:0] rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:537:3
	wire result_is_special_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:538:3
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] special_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:539:3
	wire [4:0] special_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:541:3
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:542:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:543:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:544:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:545:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:546:3
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:547:3
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:548:3
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:549:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:550:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:551:3
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:552:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) + ((NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) : 0)] mid_pipe_spec_res_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:553:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:554:3
	reg [(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_MID_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_MID_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_MID_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_MID_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] mid_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:555:3
	reg [0:NUM_MID_REGS] mid_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:556:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:557:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:559:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:562:3
	wire [1:1] sv2v_tmp_56A72;
	assign sv2v_tmp_56A72 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_56A72;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:563:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_8565A;
	assign sv2v_tmp_8565A = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_8565A;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:564:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_F1167;
	assign sv2v_tmp_F1167 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_F1167;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:565:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_19629;
	assign sv2v_tmp_19629 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_19629;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:566:3
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_2FB0E;
	assign sv2v_tmp_2FB0E = addend_shamt + addend_normalize_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_2FB0E;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:567:3
	wire [1:1] sv2v_tmp_6F5F7;
	assign sv2v_tmp_6F5F7 = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6F5F7;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:568:3
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_74CB3;
	assign sv2v_tmp_74CB3 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_74CB3;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:569:3
	wire [1:1] sv2v_tmp_D7BD0;
	assign sv2v_tmp_D7BD0 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_D7BD0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:570:3
	wire [3:1] sv2v_tmp_2170E;
	assign sv2v_tmp_2170E = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_2170E;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:571:3
	wire [3:1] sv2v_tmp_8A4AE;
	assign sv2v_tmp_8A4AE = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_8A4AE;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:572:3
	wire [1:1] sv2v_tmp_7DEC5;
	assign sv2v_tmp_7DEC5 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_7DEC5;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:573:3
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) * 1:1] sv2v_tmp_1ADE6;
	assign sv2v_tmp_1ADE6 = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] = sv2v_tmp_1ADE6;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:574:3
	wire [5:1] sv2v_tmp_1A1E3;
	assign sv2v_tmp_1A1E3 = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_1A1E3;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:575:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_8D3DE;
	assign sv2v_tmp_8D3DE = inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	always @(*) mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_8D3DE;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:576:3
	wire [1:1] sv2v_tmp_D7646;
	assign sv2v_tmp_D7646 = inp_pipe_mask_q[NUM_INP_REGS];
	always @(*) mid_pipe_mask_q[0] = sv2v_tmp_D7646;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:577:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_E3910;
	assign sv2v_tmp_E3910 = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_E3910;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:578:3
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:580:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:583:3
	genvar _gv_i_224;
	generate
		for (_gv_i_224 = 0; _gv_i_224 < NUM_MID_REGS; _gv_i_224 = _gv_i_224 + 1) begin : gen_inside_pipeline
			localparam i = _gv_i_224;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:585:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:589:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:591:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:591:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:591:408
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:591:560
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:593:5
			assign reg_ena = (mid_pipe_ready[i] & mid_pipe_valid_q[i]) | reg_ena_i[NUM_INP_REGS + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:595:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:595:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:595:189
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:595:297
					mid_pipe_eff_sub_q[i + 1] <= (reg_ena ? mid_pipe_eff_sub_q[i] : mid_pipe_eff_sub_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:596:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:596:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:596:189
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:596:297
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:597:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:597:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:597:189
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:597:297
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:598:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:598:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:598:189
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:598:297
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:599:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:599:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:599:189
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:599:297
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= (reg_ena ? mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] : mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:600:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:600:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:600:189
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:600:297
					mid_pipe_sticky_q[i + 1] <= (reg_ena ? mid_pipe_sticky_q[i] : mid_pipe_sticky_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:601:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:601:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:601:189
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:601:297
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= (reg_ena ? mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] : mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:602:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:602:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:602:189
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:602:297
					mid_pipe_final_sign_q[i + 1] <= (reg_ena ? mid_pipe_final_sign_q[i] : mid_pipe_final_sign_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:603:89
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:603:145
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:603:201
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:603:309
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:604:101
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:604:157
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:604:213
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:604:321
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:605:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:605:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:605:189
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:605:297
					mid_pipe_res_is_spec_q[i + 1] <= (reg_ena ? mid_pipe_res_is_spec_q[i] : mid_pipe_res_is_spec_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:606:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:606:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:606:189
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:606:297
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= (reg_ena ? mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] : mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:607:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:607:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:607:189
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:607:297
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= (reg_ena ? mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5] : mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:608:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:608:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:608:199
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:608:307
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:609:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:609:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:609:189
					mid_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:609:297
					mid_pipe_mask_q[i + 1] <= (reg_ena ? mid_pipe_mask_q[i] : mid_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:610:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:610:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:610:199
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:610:307
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:613:3
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:614:3
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:615:3
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:616:3
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:617:3
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:618:3
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:619:3
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:620:3
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:621:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:622:3
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:623:3
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:624:3
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:625:3
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:630:3
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:631:3
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:632:3
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:633:3
	wire lzc_zeroes;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:635:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:636:3
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:638:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:639:3
	reg [PRECISION_BITS:0] final_mantissa;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:640:3
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:641:3
	wire sticky_after_norm;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:643:3
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:645:3
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:648:3
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:657:3
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:660:3
	always @(*) begin : norm_shift_amount
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:662:5
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:664:7
				if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:666:9
					norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:667:9
					normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
				end
				else begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:671:9
					norm_shamt = $unsigned($signed((PRECISION_BITS + 2) + exponent_product_q));
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:672:9
					normalized_exponent = 0;
				end
			end
		end
		else begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:676:7
			norm_shamt = addend_shamt_q;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:677:7
			normalized_exponent = tentative_exponent_q;
		end
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:682:3
	assign sum_shifted = sum_q << norm_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:686:3
	always @(*) begin : small_norm
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:688:5
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:689:5
		final_exponent = normalized_exponent;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:692:5
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:693:7
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:694:7
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:700:7
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:701:7
			final_exponent = normalized_exponent - 1;
		end
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:704:7
			final_exponent = 1'sb0;
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:709:3
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:714:3
	wire pre_round_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:715:3
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] pre_round_abs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:716:3
	wire [1:0] round_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:718:3
	wire of_before_round;
	wire of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:719:3
	wire uf_before_round;
	wire uf_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:721:3
	wire [(NUM_FORMATS * (SUPER_EXP_BITS + SUPER_MAN_BITS)) - 1:0] fmt_pre_round_abs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:722:3
	wire [9:0] fmt_round_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:724:3
	reg [4:0] fmt_of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:725:3
	reg [4:0] fmt_uf_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:727:3
	wire rounded_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:728:3
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] rounded_abs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:729:3
	wire result_zero;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:732:3
	assign of_before_round = final_exponent >= ((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:733:3
	assign uf_before_round = final_exponent == 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:736:3
	genvar _gv_fmt_7;
	generate
		for (_gv_fmt_7 = 0; _gv_fmt_7 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_7 = _gv_fmt_7 + 1) begin : gen_res_assemble
			localparam fmt = _gv_fmt_7;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:738:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:739:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:741:5
			wire [EXP_BITS - 1:0] pre_round_exponent;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:742:5
			wire [MAN_BITS - 1:0] pre_round_mantissa;
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:746:7
				assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : final_exponent[EXP_BITS - 1:0]);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:747:7
				assign pre_round_mantissa = (of_before_round ? {fpnew_pkg_man_bits(sv2v_cast_0BC43(_gv_fmt_7)) {1'sb1}} : final_mantissa[SUPER_MAN_BITS-:MAN_BITS]);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:749:7
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {pre_round_exponent, pre_round_mantissa};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:752:7
				assign fmt_round_sticky_bits[(fmt * 2) + 1] = final_mantissa[SUPER_MAN_BITS - MAN_BITS] | of_before_round;
				if (MAN_BITS < SUPER_MAN_BITS) begin : narrow_sticky
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:757:9
					assign fmt_round_sticky_bits[fmt * 2] = (|final_mantissa[(SUPER_MAN_BITS - MAN_BITS) - 1:0] | sticky_after_norm) | of_before_round;
				end
				else begin : normal_sticky
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:760:9
					assign fmt_round_sticky_bits[fmt * 2] = sticky_after_norm | of_before_round;
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:763:7
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {SUPER_EXP_BITS + SUPER_MAN_BITS {fpnew_pkg_DONT_CARE}};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:764:7
				assign fmt_round_sticky_bits[fmt * 2+:2] = {2 {fpnew_pkg_DONT_CARE}};
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:769:3
	assign pre_round_sign = final_sign_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:770:3
	assign pre_round_abs = fmt_pre_round_abs[dst_fmt_q2 * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:773:3
	assign round_sticky_bits = fmt_round_sticky_bits[dst_fmt_q2 * 2+:2];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:776:3
	fpnew_rounding #(.AbsWidth(SUPER_EXP_BITS + SUPER_MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:789:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:791:3
	genvar _gv_fmt_8;
	generate
		for (_gv_fmt_8 = 0; _gv_fmt_8 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_8 = _gv_fmt_8 + 1) begin : gen_sign_inject
			localparam fmt = _gv_fmt_8;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:793:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:794:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:795:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:798:7
				always @(*) begin : post_process
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:800:9
					fmt_uf_after_round[fmt] = (rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}}) || (((pre_round_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}}) && (rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == 1)) && ((round_sticky_bits != 2'b11) || (!sum_sticky_bits[(MAN_BITS * 2) + 4] && ((rnd_mode_q == 3'b000) || (rnd_mode_q == 3'b100)))));
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:803:9
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:806:9
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:807:9
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]};
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:810:7
				wire [1:1] sv2v_tmp_4A747;
				assign sv2v_tmp_4A747 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4A747;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:811:7
				wire [1:1] sv2v_tmp_90681;
				assign sv2v_tmp_90681 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_90681;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:812:7
				wire [WIDTH * 1:1] sv2v_tmp_143A7;
				assign sv2v_tmp_143A7 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_143A7;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:817:3
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:818:3
	assign of_after_round = fmt_of_after_round[dst_fmt_q2];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:824:3
	wire [WIDTH - 1:0] regular_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:825:3
	wire [4:0] regular_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:828:3
	assign regular_result = fmt_result[dst_fmt_q2 * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:829:3
	assign regular_status[4] = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:830:3
	assign regular_status[3] = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:831:3
	assign regular_status[2] = of_before_round | of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:832:3
	assign regular_status[1] = uf_after_round & regular_status[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:833:3
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:836:3
	wire [WIDTH - 1:0] result_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:837:3
	wire [4:0] status_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:840:3
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:841:3
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:847:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:848:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:849:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] out_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:850:3
	reg [0:NUM_OUT_REGS] out_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:851:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:852:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:854:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:857:3
	wire [WIDTH * 1:1] sv2v_tmp_1212D;
	assign sv2v_tmp_1212D = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_1212D;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:858:3
	wire [5:1] sv2v_tmp_F691B;
	assign sv2v_tmp_F691B = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_F691B;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:859:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_D7037;
	assign sv2v_tmp_D7037 = mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_D7037;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:860:3
	wire [1:1] sv2v_tmp_DB780;
	assign sv2v_tmp_DB780 = mid_pipe_mask_q[NUM_MID_REGS];
	always @(*) out_pipe_mask_q[0] = sv2v_tmp_DB780;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:861:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_E6477;
	assign sv2v_tmp_E6477 = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_E6477;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:862:3
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:864:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:866:3
	genvar _gv_i_225;
	generate
		for (_gv_i_225 = 0; _gv_i_225 < NUM_OUT_REGS; _gv_i_225 = _gv_i_225 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_225;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:868:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:872:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:874:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:874:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:874:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:874:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:876:5
			assign reg_ena = (out_pipe_ready[i] & out_pipe_valid_q[i]) | reg_ena_i[(NUM_INP_REGS + NUM_MID_REGS) + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:878:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:878:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:878:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:878:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:879:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:879:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:879:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:879:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:880:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:880:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:880:189
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:880:297
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:881:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:881:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:881:179
					out_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:881:287
					out_pipe_mask_q[i + 1] <= (reg_ena ? out_pipe_mask_q[i] : out_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:882:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:882:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:882:189
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:882:297
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:885:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:887:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:888:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:889:3
	assign extension_bit_o = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:890:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:891:3
	assign mask_o = out_pipe_mask_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:892:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:893:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma_multi.sv:894:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_rounding (
	abs_value_i,
	sign_i,
	round_sticky_bits_i,
	rnd_mode_i,
	effective_subtraction_i,
	abs_rounded_o,
	sign_o,
	exact_zero_o
);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:17:13
	parameter [31:0] AbsWidth = 2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:20:3
	input wire [AbsWidth - 1:0] abs_value_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:21:3
	input wire sign_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:23:3
	input wire [1:0] round_sticky_bits_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:24:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:25:3
	input wire effective_subtraction_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:27:3
	output wire [AbsWidth - 1:0] abs_rounded_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:28:3
	output wire sign_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:30:3
	output wire exact_zero_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:33:3
	reg round_up;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:45:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	always @(*) begin : rounding_decision
		// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:46:5
		case (rnd_mode_i)
			3'b000:
				case (round_sticky_bits_i)
					2'b00, 2'b01:
						// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:50:18
						round_up = 1'b0;
					2'b10:
						// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:51:18
						round_up = abs_value_i[0];
					2'b11:
						// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:52:18
						round_up = 1'b1;
					default:
						// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:53:20
						round_up = fpnew_pkg_DONT_CARE;
				endcase
			3'b001:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:55:23
				round_up = 1'b0;
			3'b010:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:56:23
				round_up = (|round_sticky_bits_i ? sign_i : 1'b0);
			3'b011:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:57:23
				round_up = (|round_sticky_bits_i ? ~sign_i : 1'b0);
			3'b100:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:58:23
				round_up = round_sticky_bits_i[1];
			3'b101:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:59:23
				round_up = ~abs_value_i[0] & |round_sticky_bits_i;
			default:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:60:16
				round_up = fpnew_pkg_DONT_CARE;
		endcase
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:65:3
	assign abs_rounded_o = abs_value_i + round_up;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:68:3
	assign exact_zero_o = (abs_value_i == {AbsWidth {1'sb0}}) && (round_sticky_bits_i == {2 {1'sb0}});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_rounding.sv:72:3
	assign sign_o = (exact_zero_o && effective_subtraction_i ? rnd_mode_i == 3'b010 : sign_i);
endmodule
module fpnew_divsqrt_th_64_multi_5F898_8E3CD (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	dst_fmt_i,
	tag_i,
	mask_i,
	aux_i,
	vectorial_op_i,
	in_valid_i,
	in_ready_o,
	divsqrt_done_o,
	simd_synch_done_i,
	divsqrt_ready_o,
	simd_synch_rdy_i,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	mask_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o,
	reg_ena_i
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// removed localparam type TagType_TagType_TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:21:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:23:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:24:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:25:38
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:26:38
	// removed localparam type AuxType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:28:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:307:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:319:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:320:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:5
			begin : sv2v_autoblock_1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:323:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:29:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:30:14
	localparam [31:0] ExtRegEnaWidth = (NumPipeRegs == 0 ? 1 : NumPipeRegs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:32:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:33:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:35:3
	input wire [(2 * WIDTH) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:36:3
	input wire [9:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:37:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:38:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:39:3
	input wire [2:0] dst_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:40:3
	input wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:41:3
	input wire mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:42:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:43:3
	input wire vectorial_op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:45:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:46:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:47:3
	output wire divsqrt_done_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:48:3
	input wire simd_synch_done_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:49:3
	output wire divsqrt_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:50:3
	input wire simd_synch_rdy_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:51:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:53:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:54:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:55:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:56:3
	output wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:57:3
	output wire mask_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:58:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:60:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:61:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:63:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:65:3
	input wire [ExtRegEnaWidth - 1:0] reg_ena_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:72:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:77:3
	localparam NUM_OUT_REGS = ((PipeConfig == 2'd1) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:87:3
	wire [(2 * WIDTH) - 1:0] operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:88:3
	wire [2:0] rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:89:3
	wire [3:0] op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:90:3
	wire [2:0] dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:91:3
	wire in_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:94:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:95:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:96:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:97:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:98:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] inp_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:99:3
	reg [0:NUM_INP_REGS] inp_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:100:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:101:3
	reg [0:NUM_INP_REGS] inp_pipe_vec_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:102:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:104:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:107:3
	wire [2 * WIDTH:1] sv2v_tmp_2997B;
	assign sv2v_tmp_2997B = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_2997B;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:108:3
	wire [3:1] sv2v_tmp_4AE25;
	assign sv2v_tmp_4AE25 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_4AE25;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:109:3
	wire [4:1] sv2v_tmp_5E107;
	assign sv2v_tmp_5E107 = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_5E107;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:110:3
	wire [3:1] sv2v_tmp_97441;
	assign sv2v_tmp_97441 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_97441;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:111:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_94CC2;
	assign sv2v_tmp_94CC2 = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_94CC2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:112:3
	wire [1:1] sv2v_tmp_407DF;
	assign sv2v_tmp_407DF = mask_i;
	always @(*) inp_pipe_mask_q[0] = sv2v_tmp_407DF;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:113:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_142AF;
	assign sv2v_tmp_142AF = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_142AF;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:114:3
	wire [1:1] sv2v_tmp_EFF0C;
	assign sv2v_tmp_EFF0C = vectorial_op_i;
	always @(*) inp_pipe_vec_op_q[0] = sv2v_tmp_EFF0C;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:115:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:117:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:119:3
	genvar _gv_i_226;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] sv2v_cast_48BE4;
		input reg [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] inp;
		sv2v_cast_48BE4 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (_gv_i_226 = 0; _gv_i_226 < NUM_INP_REGS; _gv_i_226 = _gv_i_226 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_226;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:121:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:125:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:127:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:127:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:127:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:127:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:129:5
			assign reg_ena = (inp_pipe_ready[i] & inp_pipe_valid_q[i]) | reg_ena_i[i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:131:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:131:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:131:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:131:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:132:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:132:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:132:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:132:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:133:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:133:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:133:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:133:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:134:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:134:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:134:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:134:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:135:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:135:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:135:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:135:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:136:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:136:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:136:183
					inp_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:136:291
					inp_pipe_mask_q[i + 1] <= (reg_ena ? inp_pipe_mask_q[i] : inp_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:137:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:137:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:137:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:137:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:138:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:138:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:138:193
					inp_pipe_vec_op_q[i + 1] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:138:301
					inp_pipe_vec_op_q[i + 1] <= (reg_ena ? inp_pipe_vec_op_q[i] : inp_pipe_vec_op_q[i + 1]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:141:3
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:142:3
	assign rnd_mode_q = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:143:3
	assign op_q = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:144:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:145:3
	assign in_valid_q = inp_pipe_valid_q[NUM_INP_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:147:3
	wire last_inp_reg_ena;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:148:3
	generate
		if (NUM_INP_REGS >= 1) begin : gen_last_inp_reg_ena_valid
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:149:5
			assign last_inp_reg_ena = reg_ena_i[NUM_INP_REGS - 1];
		end
		else begin : gen_last_inp_reg_ena_zero
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:151:5
			assign last_inp_reg_ena = 1'b0;
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:154:3
	reg ext_op_start_q;
	// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:155:46
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:155:102
		if (!rst_ni)
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:155:158
			ext_op_start_q <= 1'b0;
		else
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:155:266
			ext_op_start_q <= last_inp_reg_ena;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:160:3
	reg [3:0] divsqrt_fmt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:163:3
	generate
		if (WIDTH == 64) begin : translate_fmt_64_bits
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:164:5
			always @(*) begin : translate_fmt
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:165:7
				case (dst_fmt_q)
					sv2v_cast_0BC43('d1):
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:166:29
						divsqrt_fmt = 4'b1000;
					sv2v_cast_0BC43('d0):
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:167:29
						divsqrt_fmt = 4'b0100;
					sv2v_cast_0BC43('d2):
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:168:29
						divsqrt_fmt = 4'b0010;
					sv2v_cast_0BC43('d4):
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:169:29
						divsqrt_fmt = 4'b0001;
					default:
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:170:29
						divsqrt_fmt = 4'b1000;
				endcase
			end
		end
		else if (WIDTH == 32) begin : translate_fmt_32_bits
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:174:5
			always @(*) begin : translate_fmt
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:175:7
				case (dst_fmt_q)
					sv2v_cast_0BC43('d0):
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:176:29
						divsqrt_fmt = 4'b0100;
					sv2v_cast_0BC43('d2):
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:177:29
						divsqrt_fmt = 4'b0010;
					sv2v_cast_0BC43('d4):
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:178:29
						divsqrt_fmt = 4'b0001;
					default:
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:179:29
						divsqrt_fmt = 4'b0100;
				endcase
			end
		end
		else if (WIDTH == 16) begin : translate_fmt_16_bits
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:183:5
			always @(*) begin : translate_fmt
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:184:7
				case (dst_fmt_q)
					sv2v_cast_0BC43('d2):
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:185:29
						divsqrt_fmt = 4'b0010;
					sv2v_cast_0BC43('d4):
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:186:29
						divsqrt_fmt = 4'b0001;
					default:
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:187:29
						divsqrt_fmt = 4'b0010;
				endcase
			end
		end
		else begin : genblk3
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:191:5
			$fatal(1, "DivSqrt THMULTI: Unsupported WIDTH (the supported width are 64, 32, 16)");
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:198:3
	reg in_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:199:3
	wire div_valid;
	wire sqrt_valid;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:200:3
	wire unit_ready;
	wire unit_done;
	reg unit_done_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:201:3
	wire op_starting;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:202:3
	reg out_valid;
	wire out_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:203:3
	reg unit_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:204:3
	wire simd_synch_done;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:206:3
	// removed localparam type fsm_state_e
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:207:3
	reg [1:0] state_q;
	reg [1:0] state_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:210:3
	assign div_valid = (((in_valid_q & in_ready) & ~flush_i) | ext_op_start_q) & (op_q == sv2v_cast_A53F3(4));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:211:3
	assign sqrt_valid = (((in_valid_q & in_ready) & ~flush_i) | ext_op_start_q) & (op_q != sv2v_cast_A53F3(4));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:212:3
	assign op_starting = div_valid | sqrt_valid;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:216:3
	reg [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] result_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:217:3
	reg result_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:218:3
	reg [AuxType_AUX_BITS - 1:0] result_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:219:3
	reg result_vec_op_q;
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:222:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:222:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:222:182
			result_tag_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:222:290
			result_tag_q <= (op_starting ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : result_tag_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:223:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:223:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:223:182
			result_mask_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:223:290
			result_mask_q <= (op_starting ? inp_pipe_mask_q[NUM_INP_REGS] : result_mask_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:224:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:224:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:224:182
			result_aux_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:224:290
			result_aux_q <= (op_starting ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : result_aux_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:225:73
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:225:129
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:225:185
			result_vec_op_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:225:293
			result_vec_op_q <= (op_starting ? inp_pipe_vec_op_q[NUM_INP_REGS] : result_vec_op_q);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:228:3
	assign simd_synch_done = simd_synch_done_i || ~result_vec_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:233:3
	wire unit_done_clear;
	// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:234:230
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:234:308
		if (!rst_ni)
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:234:386
			unit_done_q <= 1'b0;
		else
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:234:538
			unit_done_q <= (unit_done_clear ? 1'b0 : (unit_done ? unit_done : unit_done_q));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:235:3
	assign unit_done_clear = simd_synch_done | last_inp_reg_ena;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:237:3
	assign divsqrt_done_o = (unit_done_q | unit_done) & result_vec_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:241:3
	assign divsqrt_ready_o = in_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:243:3
	assign inp_pipe_ready[NUM_INP_REGS] = (result_vec_op_q ? simd_synch_rdy_i : in_ready);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:246:3
	always @(*) begin : flag_fsm
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:248:5
		in_ready = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:249:5
		out_valid = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:250:5
		unit_busy = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:251:5
		state_d = state_q;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:253:5
		case (state_q)
			2'd0: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:256:9
				in_ready = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:257:9
				if (in_valid_q && unit_ready)
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:258:11
					state_d = 2'd1;
			end
			2'd1: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:263:9
				unit_busy = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:265:9
				if (simd_synch_done_i || (~result_vec_op_q && unit_done)) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:266:11
					out_valid = 1'b1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:268:11
					if (out_ready) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:269:13
						state_d = 2'd0;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:270:13
						in_ready = 1'b1;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:271:13
						if (in_valid_q && unit_ready)
							// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:272:15
							state_d = 2'd1;
					end
					else
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:276:13
						state_d = 2'd2;
				end
			end
			2'd2: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:282:9
				unit_busy = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:283:9
				out_valid = 1'b1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:285:9
				if (out_ready) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:286:11
					state_d = 2'd0;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:287:11
					if (in_valid_q && unit_ready) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:288:13
						in_ready = 1'b1;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:289:13
						state_d = 2'd1;
					end
				end
			end
			default:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:294:16
				state_d = 2'd0;
		endcase
		if (flush_i) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:299:7
			unit_busy = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:300:7
			out_valid = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:301:7
			state_d = 2'd0;
		end
	end
	// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:306:30
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:306:86
		if (!rst_ni)
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:306:142
			state_q <= 2'd0;
		else
			// Trace: macro expansion of FF at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:306:250
			state_q <= state_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:311:3
	wire [63:0] unit_result;
	reg [63:0] held_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:312:3
	wire [4:0] unit_status;
	reg [4:0] held_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:313:3
	wire hold_en;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:315:3
	wire vfdsu_dp_fdiv_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:318:3
	reg [2:0] rm_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:319:3
	reg [3:0] divsqrt_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:320:3
	reg [3:0] divsqrt_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:321:3
	wire div_op;
	wire sqrt_op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:322:3
	reg [WIDTH - 1:0] srcf0_q;
	reg [WIDTH - 1:0] srcf1_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:323:3
	reg [63:0] srcf0;
	reg [63:0] srcf1;
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:326:53
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:326:109
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:326:165
			rm_q <= 3'b000;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:326:273
			rm_q <= (op_starting ? rnd_mode_q : rm_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:327:51
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:327:107
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:327:163
			divsqrt_fmt_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:327:271
			divsqrt_fmt_q <= (op_starting ? divsqrt_fmt : divsqrt_fmt_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:328:55
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:328:111
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:328:167
			divsqrt_op_q <= sv2v_cast_A53F3(4);
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:328:275
			divsqrt_op_q <= (op_starting ? op_q : divsqrt_op_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:329:47
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:329:103
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:329:159
			srcf0_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:329:267
			srcf0_q <= (op_starting ? operands_q[0+:WIDTH] : srcf0_q);
	// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:330:47
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:330:103
		if (!rst_ni)
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:330:159
			srcf1_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:330:267
			srcf1_q <= (op_starting ? operands_q[WIDTH+:WIDTH] : srcf1_q);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:333:3
	generate
		if (WIDTH == 64) begin : gen_fmt_64_bits
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:334:5
			always @(*) begin : NaN_box_inputs
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:335:7
				if (divsqrt_fmt_q == 4'b1000) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:336:9
					srcf0[63:0] = srcf0_q[63:0];
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:337:9
					srcf1[63:0] = srcf1_q[63:0];
				end
				else if (divsqrt_fmt_q == 4'b0100) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:339:9
					srcf0[63:32] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:340:9
					srcf1[63:32] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:341:9
					srcf0[31:0] = srcf0_q[31:0];
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:342:9
					srcf1[31:0] = srcf1_q[31:0];
				end
				else if ((divsqrt_fmt_q == 4'b0010) || (divsqrt_fmt_q == 4'b0001)) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:344:9
					srcf0[63:16] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:345:9
					srcf1[63:16] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:346:9
					srcf0[15:0] = srcf0_q[15:0];
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:347:9
					srcf1[15:0] = srcf1_q[15:0];
				end
				else begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:349:9
					srcf0[63:0] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:350:9
					srcf1[63:0] = 1'sb1;
				end
			end
		end
		else if (WIDTH == 32) begin : gen_fmt_32_bits
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:354:5
			always @(*) begin : NaN_box_inputs
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:355:7
				if (divsqrt_fmt_q == 4'b0100) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:356:9
					srcf0[63:32] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:357:9
					srcf1[63:32] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:358:9
					srcf0[31:0] = srcf0_q[31:0];
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:359:9
					srcf1[31:0] = srcf1_q[31:0];
				end
				else if ((divsqrt_fmt_q == 4'b0010) || (divsqrt_fmt_q == 4'b0001)) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:361:9
					srcf0[63:16] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:362:9
					srcf1[63:16] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:363:9
					srcf0[15:0] = srcf0_q[15:0];
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:364:9
					srcf1[15:0] = srcf1_q[15:0];
				end
				else begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:366:9
					srcf0[63:0] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:367:9
					srcf1[63:0] = 1'sb1;
				end
			end
		end
		else if (WIDTH == 16) begin : gen_fmt_16_bits
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:371:5
			always @(*) begin : NaN_box_inputs
				// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:372:7
				if ((divsqrt_fmt_q == 4'b0010) || (divsqrt_fmt_q == 4'b0001)) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:373:9
					srcf0[63:16] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:374:9
					srcf1[63:16] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:375:9
					srcf0[15:0] = srcf0_q[15:0];
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:376:9
					srcf1[15:0] = srcf1_q[15:0];
				end
				else begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:378:9
					srcf0[63:0] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:379:9
					srcf1[63:0] = 1'sb1;
				end
			end
		end
		else begin : genblk4
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:383:5
			$fatal(1, "DivSqrt THMULTI: Unsupported WIDTH (the supported width are 64, 32, 16)");
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:386:3
	assign div_op = (divsqrt_op_q == sv2v_cast_A53F3(4) ? 1'b1 : 1'b0);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:387:3
	assign sqrt_op = (divsqrt_op_q != sv2v_cast_A53F3(4) ? 1'b1 : 1'b0);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:390:3
	reg func_sel;
	// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:391:217
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:391:295
		if (!rst_ni)
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:391:373
			func_sel <= 1'b0;
		else
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:391:525
			func_sel <= (func_sel ? 1'b0 : (op_starting ? 1'b1 : func_sel));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:394:3
	reg op_sel;
	// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:395:210
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:395:288
		if (!rst_ni)
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:395:366
			op_sel <= 1'b0;
		else
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:395:518
			op_sel <= (op_sel ? 1'b0 : (func_sel ? 1'b1 : op_sel));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:397:3
	ct_vfdsu_top i_ct_vfdsu_top(
		.cp0_vfpu_icg_en(1'b0),
		.cp0_yy_clk_en(1'b1),
		.cpurst_b(rst_ni),
		.dp_vfdsu_ex1_pipex_dst_ereg(1'sb0),
		.dp_vfdsu_ex1_pipex_dst_vreg(1'sb0),
		.dp_vfdsu_ex1_pipex_iid(1'sb0),
		.dp_vfdsu_ex1_pipex_imm0(3'b111),
		.dp_vfdsu_ex1_pipex_sel(op_sel),
		.dp_vfdsu_ex1_pipex_srcf0(srcf0),
		.dp_vfdsu_ex1_pipex_srcf1(srcf1),
		.dp_vfdsu_fdiv_gateclk_issue(1'b1),
		.dp_vfdsu_idu_fdiv_issue(op_starting),
		.forever_cpuclk(clk_i),
		.idu_vfpu_rf_pipex_func({3'b000, divsqrt_fmt_q, 11'b00000000000, sqrt_op, div_op}),
		.idu_vfpu_rf_pipex_gateclk_sel(func_sel),
		.pad_yy_icg_scan_en(1'b0),
		.rtu_yy_xx_flush(flush_i | last_inp_reg_ena),
		.vfpu_yy_xx_dqnan(1'b0),
		.vfpu_yy_xx_rm(rm_q),
		.pipex_dp_vfdsu_ereg(),
		.pipex_dp_vfdsu_ereg_data(unit_status),
		.pipex_dp_vfdsu_freg_data(unit_result),
		.pipex_dp_vfdsu_inst_vld(unit_done),
		.pipex_dp_vfdsu_vreg(),
		.vfdsu_dp_fdiv_busy(vfdsu_dp_fdiv_busy),
		.vfdsu_dp_inst_wb_req(),
		.vfdsu_ifu_debug_ex2_wait(),
		.vfdsu_ifu_debug_idle(),
		.vfdsu_ifu_debug_pipe_busy()
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:429:3
	assign unit_ready = !vfdsu_dp_fdiv_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:433:3
	assign hold_en = (unit_done & (~simd_synch_done_i | ~out_ready)) & ~(~result_vec_op_q & out_ready);
	// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:435:50
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:435:92
		held_result_q <= (hold_en ? unit_result : held_result_q);
	// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:436:50
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:436:92
		held_status_q <= (hold_en ? unit_status : held_status_q);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:441:3
	wire [WIDTH - 1:0] result_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:442:3
	wire [4:0] status_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:444:3
	assign result_d[WIDTH - 1:0] = (unit_done_q ? held_result_q[WIDTH - 1:0] : unit_result[WIDTH - 1:0]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:445:3
	assign status_d = (unit_done_q ? held_status_q : unit_status);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:451:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:452:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:453:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] out_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:454:3
	reg [0:NUM_OUT_REGS] out_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:455:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:456:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:458:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:461:3
	wire [WIDTH * 1:1] sv2v_tmp_E054D;
	assign sv2v_tmp_E054D = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_E054D;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:462:3
	wire [5:1] sv2v_tmp_C248B;
	assign sv2v_tmp_C248B = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_C248B;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:463:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_815FC;
	assign sv2v_tmp_815FC = result_tag_q;
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_815FC;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:464:3
	wire [1:1] sv2v_tmp_11413;
	assign sv2v_tmp_11413 = result_mask_q;
	always @(*) out_pipe_mask_q[0] = sv2v_tmp_11413;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:465:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_2F6CD;
	assign sv2v_tmp_2F6CD = result_aux_q;
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_2F6CD;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:466:3
	wire [1:1] sv2v_tmp_D06FD;
	assign sv2v_tmp_D06FD = out_valid;
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_D06FD;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:468:3
	assign out_ready = out_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:470:3
	genvar _gv_i_227;
	generate
		for (_gv_i_227 = 0; _gv_i_227 < NUM_OUT_REGS; _gv_i_227 = _gv_i_227 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_227;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:472:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:476:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:478:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:478:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:478:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:478:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:480:5
			assign reg_ena = (out_pipe_ready[i] & out_pipe_valid_q[i]) | reg_ena_i[NUM_INP_REGS + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:482:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:482:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:482:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:482:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:483:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:483:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:483:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:483:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:484:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:484:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:484:189
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:484:297
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:485:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:485:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:485:179
					out_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:485:287
					out_pipe_mask_q[i + 1] <= (reg_ena ? out_pipe_mask_q[i] : out_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:486:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:486:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:486:189
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:486:297
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:489:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:491:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:492:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:493:3
	assign extension_bit_o = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:494:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:495:3
	assign mask_o = out_pipe_mask_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:496:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:497:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_divsqrt_th_64_multi.sv:498:3
	assign busy_o = |{inp_pipe_valid_q, unit_busy, out_pipe_valid_q};
endmodule
module fpnew_opgroup_fmt_slice_F5668_FC739 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	vectorial_op_i,
	tag_i,
	simd_mask_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o,
	reg_ena_i
);
	// removed localparam type TagType_TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:17:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:18:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:20:13
	parameter [31:0] Width = 32;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:21:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:22:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:23:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:24:13
	parameter [0:0] ExtRegEna = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:25:38
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:26:13
	parameter [31:0] TrueSIMDClass = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:28:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:389:48
		input reg [1:0] grp;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:390:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:29:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic [31:0] fpnew_pkg_num_lanes;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:400:45
		input reg [31:0] width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:400:65
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:400:82
		input reg vec;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:401:5
		fpnew_pkg_num_lanes = (vec ? width / fpnew_pkg_fp_width(fmt) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_num_lanes(Width, FpFormat, EnableVectors);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:30:27
	// removed localparam type MaskType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:31:14
	localparam [31:0] ExtRegEnaWidth = (NumPipeRegs == 0 ? 1 : NumPipeRegs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:33:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:34:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:36:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:37:3
	input wire [NUM_OPERANDS - 1:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:38:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:39:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:40:3
	input wire op_mod_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:41:3
	input wire vectorial_op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:42:3
	input wire [TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:43:3
	input wire [NUM_LANES - 1:0] simd_mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:45:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:46:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:47:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:49:3
	output wire [Width - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:50:3
	// removed localparam type fpnew_pkg_status_t
	output reg [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:51:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:52:3
	output wire [TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:54:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:55:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:57:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:59:3
	input wire [ExtRegEnaWidth - 1:0] reg_ena_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:62:3
	localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:63:3
	localparam [31:0] SIMD_WIDTH = $unsigned(Width / NUM_LANES);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:66:3
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:67:3
	wire vectorial_op;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:69:3
	wire [(NUM_LANES * FP_WIDTH) - 1:0] slice_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:70:3
	wire [Width - 1:0] slice_regular_result;
	wire [Width - 1:0] slice_class_result;
	wire [Width - 1:0] slice_vec_class_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:72:3
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:73:3
	wire [NUM_LANES - 1:0] lane_ext_bit;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:74:3
	// removed localparam type fpnew_pkg_classmask_e
	wire [(NUM_LANES * 10) - 1:0] lane_class_mask;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:75:3
	wire [((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? (NUM_LANES * (TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : (NUM_LANES * (1 - (TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TAG_WIDTH - 1)):((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0)] lane_tags;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:76:3
	wire [NUM_LANES - 1:0] lane_masks;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:77:3
	wire [NUM_LANES - 1:0] lane_vectorial;
	wire [NUM_LANES - 1:0] lane_busy;
	wire [NUM_LANES - 1:0] lane_is_class;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:79:3
	wire result_is_vector;
	wire result_is_class;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:84:3
	assign in_ready_o = lane_in_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:85:3
	assign vectorial_op = vectorial_op_i & EnableVectors;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:90:3
	genvar _gv_lane_2;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_lane_2 = 0; _gv_lane_2 < sv2v_cast_32_signed(NUM_LANES); _gv_lane_2 = _gv_lane_2 + 1) begin : gen_num_lanes
			localparam lane = _gv_lane_2;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:91:5
			wire [FP_WIDTH - 1:0] local_result;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:92:5
			wire local_sign;
			if ((lane == 0) || EnableVectors) begin : active_lane
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:96:7
				wire in_valid;
				wire out_valid;
				wire out_ready;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:98:7
				reg [(NUM_OPERANDS * FP_WIDTH) - 1:0] local_operands;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:99:7
				wire [FP_WIDTH - 1:0] op_result;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:100:7
				wire [4:0] op_status;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:102:7
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:104:7
				always @(*) begin : prepare_input
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:105:9
					begin : sv2v_autoblock_1
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:105:14
						reg signed [31:0] i;
						// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:105:14
						for (i = 0; i < sv2v_cast_32_signed(NUM_OPERANDS); i = i + 1)
							begin
								// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:106:11
								local_operands[i * FP_WIDTH+:FP_WIDTH] = operands_i[(i * Width) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (($unsigned(lane) + 1) * FP_WIDTH) - 1 : (((($unsigned(lane) + 1) * FP_WIDTH) - 1) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:(((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)];
							end
					end
				end
				if (OpGroup == 2'd0) begin : lane_instance
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:112:9
					fpnew_fma_7C8F3_7759B #(
						.TagType_TagType_TagType_TagType_TAG_WIDTH(TagType_TagType_TagType_TAG_WIDTH),
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fma(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.mask_i(simd_mask_i[lane]),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + (lane * ((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))]),
						.mask_o(lane_masks[lane]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane]),
						.reg_ena_i(reg_ena_i)
					);
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:143:9
					assign lane_is_class[lane] = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:144:9
					assign lane_class_mask[lane * 10+:10] = 10'b0000000001;
				end
				else if (OpGroup == 2'd1) begin
					;
				end
				else if (OpGroup == 2'd2) begin : lane_instance
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:177:9
					fpnew_noncomp_59FAB_0570D #(
						.TagType_TagType_TagType_TagType_TAG_WIDTH(TagType_TagType_TagType_TAG_WIDTH),
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_noncomp(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.mask_i(simd_mask_i[lane]),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.class_mask_o(lane_class_mask[lane * 10+:10]),
						.is_class_o(lane_is_class[lane]),
						.tag_o(lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + (lane * ((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))]),
						.mask_o(lane_masks[lane]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane]),
						.reg_ena_i(reg_ena_i)
					);
				end
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:213:7
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:214:7
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:217:7
				assign local_result = (lane_out_valid[lane] | ExtRegEna ? op_result : {FP_WIDTH {lane_ext_bit[0]}});
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:218:7
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] | ExtRegEna ? op_status : {5 {1'sb0}});
			end
			else begin : genblk1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:222:7
				assign lane_out_valid[lane] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:223:7
				assign lane_in_ready[lane] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:224:7
				assign local_result = {FP_WIDTH {lane_ext_bit[0]}};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:225:7
				assign lane_status[lane * 5+:5] = 1'sb0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:226:7
				assign lane_busy[lane] = 1'b0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:227:7
				assign lane_is_class[lane] = 1'b0;
			end
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:231:5
			assign slice_result[(($unsigned(lane) + 1) * FP_WIDTH) - 1:$unsigned(lane) * FP_WIDTH] = local_result;
			if (TrueSIMDClass && (SIMD_WIDTH >= 10)) begin : vectorial_true_class
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:235:7
				assign slice_vec_class_result[lane * SIMD_WIDTH+:10] = lane_class_mask[lane * 10+:10];
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:236:7
				assign slice_vec_class_result[((lane + 1) * SIMD_WIDTH) - 1-:SIMD_WIDTH - 10] = 1'sb0;
			end
			else if (((lane + 1) * 8) <= Width) begin : vectorial_class
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:238:7
				assign local_sign = (((lane_class_mask[lane * 10+:10] == 10'b0000000001) || (lane_class_mask[lane * 10+:10] == 10'b0000000010)) || (lane_class_mask[lane * 10+:10] == 10'b0000000100)) || (lane_class_mask[lane * 10+:10] == 10'b0000001000);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:243:7
				assign slice_vec_class_result[((lane + 1) * 8) - 1:lane * 8] = {local_sign, ~local_sign, lane_class_mask[lane * 10+:10] == 10'b1000000000, lane_class_mask[lane * 10+:10] == 10'b0100000000, (lane_class_mask[lane * 10+:10] == 10'b0000010000) || (lane_class_mask[lane * 10+:10] == 10'b0000001000), (lane_class_mask[lane * 10+:10] == 10'b0000100000) || (lane_class_mask[lane * 10+:10] == 10'b0000000100), (lane_class_mask[lane * 10+:10] == 10'b0001000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000010), (lane_class_mask[lane * 10+:10] == 10'b0010000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000001)};
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:263:3
	assign result_is_vector = lane_vectorial[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:264:3
	assign result_is_class = lane_is_class[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:266:3
	assign slice_regular_result = $signed({extension_bit_o, slice_result});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:268:3
	localparam [31:0] CLASS_VEC_BITS = ((NUM_LANES * 8) > Width ? 8 * (Width / 8) : NUM_LANES * 8);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:271:3
	generate
		if (!(TrueSIMDClass && (SIMD_WIDTH >= 10))) begin : genblk2
			if (CLASS_VEC_BITS < Width) begin : pad_vectorial_class
				// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:273:7
				assign slice_vec_class_result[Width - 1:CLASS_VEC_BITS] = 1'sb0;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:279:3
	assign slice_class_result = (result_is_vector ? slice_vec_class_result : lane_class_mask[0+:10]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:282:3
	assign result_o = (result_is_class ? slice_class_result : slice_regular_result);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:284:3
	assign extension_bit_o = lane_ext_bit[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:285:3
	assign tag_o = lane_tags[((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TAG_WIDTH + 0) + 0+:((TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:286:3
	assign busy_o = |lane_busy;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:287:3
	assign out_valid_o = lane_out_valid[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:291:3
	always @(*) begin : output_processing
		// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:293:5
		reg [4:0] temp_status;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:294:5
		temp_status = 1'sb0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:295:5
		begin : sv2v_autoblock_2
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:295:10
			reg signed [31:0] i;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:295:10
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:296:7
					temp_status = temp_status | (lane_status[i * 5+:5] & {5 {lane_masks[i]}});
				end
		end
		// Trace: /vortex/third_party/cvfpu/src/fpnew_opgroup_fmt_slice.sv:297:5
		status_o = temp_status;
	end
endmodule
module fpnew_cast_multi_ACFE7_57164 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	tag_i,
	mask_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	mask_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o,
	reg_ena_i
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// removed localparam type TagType_TagType_TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:19:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:20:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtConfig = 1'sb1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:22:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:23:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:24:38
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:25:38
	// removed localparam type AuxType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:27:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:307:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:319:48
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:320:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:5
			begin : sv2v_autoblock_1
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				reg [31:0] i;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:321:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:323:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:88:45
		input reg [1:0] ifmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:89:5
		case (ifmt)
			sv2v_cast_87CC5(0): fpnew_pkg_int_width = 8;
			sv2v_cast_87CC5(1): fpnew_pkg_int_width = 16;
			sv2v_cast_87CC5(2): fpnew_pkg_int_width = 32;
			sv2v_cast_87CC5(3): fpnew_pkg_int_width = 64;
			default: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:96:9
				$fatal(1, "Invalid INT format supplied");
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:100:9
				fpnew_pkg_int_width = sv2v_cast_87CC5(0);
			end
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:366:49
		input reg [0:3] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:367:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:368:5
			begin : sv2v_autoblock_2
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:368:10
				reg signed [31:0] ifmt;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:368:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:369:7
						if (cfg[ifmt])
							// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:369:22
							res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)));
					end
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_maximum(fpnew_pkg_max_fp_width(FpFmtConfig), fpnew_pkg_max_int_width(IntFmtConfig));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:29:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:30:14
	localparam [31:0] ExtRegEnaWidth = (NumPipeRegs == 0 ? 1 : NumPipeRegs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:32:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:33:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:35:3
	input wire [WIDTH - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:36:3
	input wire [4:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:37:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:38:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:39:3
	input wire op_mod_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:40:3
	input wire [2:0] src_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:41:3
	input wire [2:0] dst_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:42:3
	input wire [1:0] int_fmt_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:43:3
	input wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:44:3
	input wire mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:45:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:47:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:48:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:49:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:51:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:52:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:53:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:54:3
	output wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:55:3
	output wire mask_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:56:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:58:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:59:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:61:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:63:3
	input wire [ExtRegEnaWidth - 1:0] reg_ena_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:69:3
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:70:3
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:72:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:337:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:338:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:342:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:343:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:351:49
		input reg [0:4] cfg;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:352:5
		reg [63:0] res;
		begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:353:5
			res = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:354:5
			begin : sv2v_autoblock_3
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:354:10
				reg [31:0] fmt;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:354:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:356:9
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt))));
						// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:357:9
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:74:3
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:75:3
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:76:3
	localparam [31:0] SUPER_BIAS = (2 ** (SUPER_EXP_BITS - 1)) - 1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:79:3
	localparam [31:0] INT_MAN_WIDTH = fpnew_pkg_maximum(SUPER_MAN_BITS + 1, MAX_INT_WIDTH);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:81:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(INT_MAN_WIDTH);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:84:3
	localparam [31:0] INT_EXP_WIDTH = fpnew_pkg_maximum($clog2(MAX_INT_WIDTH), fpnew_pkg_maximum(SUPER_EXP_BITS, $clog2(SUPER_BIAS + SUPER_MAN_BITS))) + 1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:87:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:92:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:97:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:107:3
	wire [WIDTH - 1:0] operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:108:3
	wire [4:0] is_boxed_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:109:3
	wire op_mod_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:110:3
	wire [2:0] src_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:111:3
	wire [2:0] dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:112:3
	wire [1:0] int_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:115:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * WIDTH) + ((NUM_INP_REGS * WIDTH) - 1) : ((NUM_INP_REGS + 1) * WIDTH) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * WIDTH : 0)] inp_pipe_operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:116:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)] inp_pipe_is_boxed_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:117:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:118:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:119:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:120:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:121:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:122:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] inp_pipe_int_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:123:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] inp_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:124:3
	reg [0:NUM_INP_REGS] inp_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:125:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:126:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:128:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:131:3
	wire [WIDTH * 1:1] sv2v_tmp_6E45B;
	assign sv2v_tmp_6E45B = operands_i;
	always @(*) inp_pipe_operands_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * WIDTH+:WIDTH] = sv2v_tmp_6E45B;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:132:3
	wire [5:1] sv2v_tmp_C47E1;
	assign sv2v_tmp_C47E1 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS] = sv2v_tmp_C47E1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:133:3
	wire [3:1] sv2v_tmp_45ED9;
	assign sv2v_tmp_45ED9 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_45ED9;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:134:3
	wire [4:1] sv2v_tmp_AD1FB;
	assign sv2v_tmp_AD1FB = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_AD1FB;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:135:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:136:3
	wire [3:1] sv2v_tmp_CB295;
	assign sv2v_tmp_CB295 = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_CB295;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:137:3
	wire [3:1] sv2v_tmp_6AF63;
	assign sv2v_tmp_6AF63 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_6AF63;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:138:3
	wire [2:1] sv2v_tmp_CA55F;
	assign sv2v_tmp_CA55F = int_fmt_i;
	always @(*) inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_CA55F;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:139:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_C893E;
	assign sv2v_tmp_C893E = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_C893E;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:140:3
	wire [1:1] sv2v_tmp_407DF;
	assign sv2v_tmp_407DF = mask_i;
	always @(*) inp_pipe_mask_q[0] = sv2v_tmp_407DF;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:141:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_73173;
	assign sv2v_tmp_73173 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_73173;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:142:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:144:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:146:3
	genvar _gv_i_228;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] sv2v_cast_48BE4;
		input reg [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] inp;
		sv2v_cast_48BE4 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (_gv_i_228 = 0; _gv_i_228 < NUM_INP_REGS; _gv_i_228 = _gv_i_228 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_228;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:148:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:152:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:154:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:154:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:154:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:154:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:156:5
			assign reg_ena = (inp_pipe_ready[i] & inp_pipe_valid_q[i]) | reg_ena_i[i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:158:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:158:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:158:183
					inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:158:291
					inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * WIDTH+:WIDTH] : inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:159:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:159:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:159:183
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:159:291
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS+:NUM_FORMATS] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:160:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:160:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:160:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:160:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:161:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:161:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:161:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:161:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:162:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:162:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:162:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:162:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:163:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:163:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:163:207
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:163:315
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:164:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:164:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:164:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:164:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:165:96
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:165:152
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:165:208
					inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_87CC5(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:165:316
					inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= (reg_ena ? inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] : inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:166:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:166:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:166:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:166:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:167:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:167:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:167:183
					inp_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:167:291
					inp_pipe_mask_q[i + 1] <= (reg_ena ? inp_pipe_mask_q[i] : inp_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:168:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:168:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:168:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:168:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:171:3
	assign operands_q = inp_pipe_operands_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:172:3
	assign is_boxed_q = inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:173:3
	assign op_mod_q = inp_pipe_op_mod_q[NUM_INP_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:174:3
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:175:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:176:3
	assign int_fmt_q = inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:181:3
	wire src_is_int;
	wire dst_is_int;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:183:3
	assign src_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(12);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:184:3
	assign dst_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(11);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:186:3
	wire [INT_MAN_WIDTH - 1:0] encoded_mant;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:188:3
	wire [4:0] fmt_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:189:3
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_exponent;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:190:3
	wire [(NUM_FORMATS * INT_MAN_WIDTH) - 1:0] fmt_mantissa;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:191:3
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_shift_compensation;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:193:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [39:0] info;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:195:3
	reg [(NUM_INT_FORMATS * INT_MAN_WIDTH) - 1:0] ifmt_input_val;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:196:3
	wire int_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:197:3
	wire [INT_MAN_WIDTH - 1:0] int_value;
	wire [INT_MAN_WIDTH - 1:0] int_mantissa;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:200:3
	genvar _gv_fmt_9;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic signed [0:0] sv2v_cast_1_signed;
		input reg signed [0:0] inp;
		sv2v_cast_1_signed = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_fmt_9 = 0; _gv_fmt_9 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_9 = _gv_fmt_9 + 1) begin : fmt_init_inputs
			localparam fmt = _gv_fmt_9;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:202:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:203:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:204:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:207:7
				localparam [2:0] FpFormat = sv2v_cast_0BC43(fmt);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:210:7
				fpnew_classifier #(
					.FpFormat(FpFormat),
					.NumOperands(1)
				) i_fpnew_classifier(
					.operands_i(operands_q[FP_WIDTH - 1:0]),
					.is_boxed_i(is_boxed_q[fmt]),
					.info_o(info[fmt * 8+:8])
				);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:219:7
				assign fmt_sign[fmt] = operands_q[FP_WIDTH - 1];
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:220:7
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed({1'b0, operands_q[MAN_BITS+:EXP_BITS]});
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:221:7
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {info[(fmt * 8) + 7], operands_q[MAN_BITS - 1:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:223:7
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed((INT_MAN_WIDTH - 1) - MAN_BITS);
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:225:7
				assign info[fmt * 8+:8] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:226:7
				assign fmt_sign[fmt] = fpnew_pkg_DONT_CARE;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:227:7
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:228:7
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:229:7
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:234:3
	genvar _gv_ifmt_3;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	generate
		for (_gv_ifmt_3 = 0; _gv_ifmt_3 < sv2v_cast_32_signed(NUM_INT_FORMATS); _gv_ifmt_3 = _gv_ifmt_3 + 1) begin : gen_sign_extend_int
			localparam ifmt = _gv_ifmt_3;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:236:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:239:7
				always @(*) begin : sign_ext_input
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:241:9
					ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {sv2v_cast_1(operands_q[INT_WIDTH - 1] & ~op_mod_q)}};
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:242:9
					ifmt_input_val[(ifmt * INT_MAN_WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = operands_q[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:245:7
				wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_5B946;
				assign sv2v_tmp_5B946 = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_5B946;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:250:3
	assign int_value = ifmt_input_val[int_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:251:3
	assign int_sign = int_value[INT_MAN_WIDTH - 1] & ~op_mod_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:252:3
	assign int_mantissa = (int_sign ? $unsigned(-int_value) : int_value);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:255:3
	assign encoded_mant = (src_is_int ? int_mantissa : fmt_mantissa[src_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:260:3
	wire signed [INT_EXP_WIDTH - 1:0] src_bias;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:261:3
	wire signed [INT_EXP_WIDTH - 1:0] src_exp;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:262:3
	wire signed [INT_EXP_WIDTH - 1:0] src_subnormal;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:263:3
	wire signed [INT_EXP_WIDTH - 1:0] src_offset;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:265:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:347:40
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:348:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	assign src_bias = $signed(fpnew_pkg_bias(src_fmt_q));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:266:3
	assign src_exp = fmt_exponent[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:267:3
	assign src_subnormal = $signed({1'b0, info[(src_fmt_q * 8) + 6]});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:268:3
	assign src_offset = fmt_shift_compensation[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:270:3
	wire input_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:271:3
	wire signed [INT_EXP_WIDTH - 1:0] input_exp;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:272:3
	wire [INT_MAN_WIDTH - 1:0] input_mant;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:273:3
	wire mant_is_zero;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:275:3
	wire signed [INT_EXP_WIDTH - 1:0] fp_input_exp;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:276:3
	wire signed [INT_EXP_WIDTH - 1:0] int_input_exp;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:279:3
	wire [LZC_RESULT_WIDTH - 1:0] renorm_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:280:3
	wire [LZC_RESULT_WIDTH:0] renorm_shamt_sgn;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:283:3
	lzc #(
		.WIDTH(INT_MAN_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(encoded_mant),
		.cnt_o(renorm_shamt),
		.empty_o(mant_is_zero)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:291:3
	assign renorm_shamt_sgn = $signed({1'b0, renorm_shamt});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:294:3
	assign input_sign = (src_is_int ? int_sign : fmt_sign[src_fmt_q]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:296:3
	assign input_mant = encoded_mant << renorm_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:298:3
	assign fp_input_exp = $signed((((src_exp + src_subnormal) - src_bias) - renorm_shamt_sgn) + src_offset);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:300:3
	assign int_input_exp = $signed((INT_MAN_WIDTH - 1) - renorm_shamt_sgn);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:302:3
	assign input_exp = (src_is_int ? int_input_exp : fp_input_exp);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:304:3
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:307:3
	assign destination_exp = input_exp + $signed(fpnew_pkg_bias(dst_fmt_q));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:313:3
	wire input_sign_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:314:3
	wire signed [INT_EXP_WIDTH - 1:0] input_exp_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:315:3
	wire [INT_MAN_WIDTH - 1:0] input_mant_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:316:3
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:317:3
	wire src_is_int_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:318:3
	wire dst_is_int_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:319:3
	wire [7:0] info_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:320:3
	wire mant_is_zero_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:321:3
	wire op_mod_q2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:322:3
	wire [2:0] rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:323:3
	wire [2:0] src_fmt_q2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:324:3
	wire [2:0] dst_fmt_q2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:325:3
	wire [1:0] int_fmt_q2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:329:3
	reg [0:NUM_MID_REGS] mid_pipe_input_sign_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:330:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_input_exp_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:331:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_MAN_WIDTH) + ((NUM_MID_REGS * INT_MAN_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_MAN_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_MAN_WIDTH : 0)] mid_pipe_input_mant_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:332:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_dest_exp_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:333:3
	reg [0:NUM_MID_REGS] mid_pipe_src_is_int_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:334:3
	reg [0:NUM_MID_REGS] mid_pipe_dst_is_int_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:335:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 8) + ((NUM_MID_REGS * 8) - 1) : ((NUM_MID_REGS + 1) * 8) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 8 : 0)] mid_pipe_info_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:336:3
	reg [0:NUM_MID_REGS] mid_pipe_mant_zero_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:337:3
	reg [0:NUM_MID_REGS] mid_pipe_op_mod_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:338:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:339:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_src_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:340:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:341:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] mid_pipe_int_fmt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:342:3
	reg [(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_MID_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_MID_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_MID_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_MID_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] mid_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:343:3
	reg [0:NUM_MID_REGS] mid_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:344:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:345:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:347:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:350:3
	wire [1:1] sv2v_tmp_3DFAC;
	assign sv2v_tmp_3DFAC = input_sign;
	always @(*) mid_pipe_input_sign_q[0] = sv2v_tmp_3DFAC;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:351:3
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_9AB08;
	assign sv2v_tmp_9AB08 = input_exp;
	always @(*) mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_9AB08;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:352:3
	wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_3BE44;
	assign sv2v_tmp_3BE44 = input_mant;
	always @(*) mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_3BE44;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:353:3
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_F626F;
	assign sv2v_tmp_F626F = destination_exp;
	always @(*) mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_F626F;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:354:3
	wire [1:1] sv2v_tmp_3D9F8;
	assign sv2v_tmp_3D9F8 = src_is_int;
	always @(*) mid_pipe_src_is_int_q[0] = sv2v_tmp_3D9F8;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:355:3
	wire [1:1] sv2v_tmp_4E95C;
	assign sv2v_tmp_4E95C = dst_is_int;
	always @(*) mid_pipe_dst_is_int_q[0] = sv2v_tmp_4E95C;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:356:3
	wire [8:1] sv2v_tmp_48E57;
	assign sv2v_tmp_48E57 = info[src_fmt_q * 8+:8];
	always @(*) mid_pipe_info_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 8+:8] = sv2v_tmp_48E57;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:357:3
	wire [1:1] sv2v_tmp_4351A;
	assign sv2v_tmp_4351A = mant_is_zero;
	always @(*) mid_pipe_mant_zero_q[0] = sv2v_tmp_4351A;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:358:3
	wire [1:1] sv2v_tmp_88AB6;
	assign sv2v_tmp_88AB6 = op_mod_q;
	always @(*) mid_pipe_op_mod_q[0] = sv2v_tmp_88AB6;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:359:3
	wire [3:1] sv2v_tmp_32E16;
	assign sv2v_tmp_32E16 = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_32E16;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:360:3
	wire [3:1] sv2v_tmp_DE9EA;
	assign sv2v_tmp_DE9EA = src_fmt_q;
	always @(*) mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_DE9EA;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:361:3
	wire [3:1] sv2v_tmp_FC1E4;
	assign sv2v_tmp_FC1E4 = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_FC1E4;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:362:3
	wire [2:1] sv2v_tmp_2AE08;
	assign sv2v_tmp_2AE08 = int_fmt_q;
	always @(*) mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_2AE08;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:363:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_18044;
	assign sv2v_tmp_18044 = inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	always @(*) mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_18044;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:364:3
	wire [1:1] sv2v_tmp_D7646;
	assign sv2v_tmp_D7646 = inp_pipe_mask_q[NUM_INP_REGS];
	always @(*) mid_pipe_mask_q[0] = sv2v_tmp_D7646;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:365:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_BCA96;
	assign sv2v_tmp_BCA96 = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_BCA96;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:366:3
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:368:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:371:3
	genvar _gv_i_229;
	generate
		for (_gv_i_229 = 0; _gv_i_229 < NUM_MID_REGS; _gv_i_229 = _gv_i_229 + 1) begin : gen_inside_pipeline
			localparam i = _gv_i_229;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:373:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:377:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:379:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:379:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:379:408
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:379:560
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:381:5
			assign reg_ena = (mid_pipe_ready[i] & mid_pipe_valid_q[i]) | reg_ena_i[NUM_INP_REGS + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:383:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:383:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:383:187
					mid_pipe_input_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:383:295
					mid_pipe_input_sign_q[i + 1] <= (reg_ena ? mid_pipe_input_sign_q[i] : mid_pipe_input_sign_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:384:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:384:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:384:187
					mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:384:295
					mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= (reg_ena ? mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH] : mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:385:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:385:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:385:187
					mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:385:295
					mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= (reg_ena ? mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_MAN_WIDTH+:INT_MAN_WIDTH] : mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:386:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:386:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:386:187
					mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:386:295
					mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= (reg_ena ? mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH] : mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:387:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:387:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:387:187
					mid_pipe_src_is_int_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:387:295
					mid_pipe_src_is_int_q[i + 1] <= (reg_ena ? mid_pipe_src_is_int_q[i] : mid_pipe_src_is_int_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:388:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:388:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:388:187
					mid_pipe_dst_is_int_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:388:295
					mid_pipe_dst_is_int_q[i + 1] <= (reg_ena ? mid_pipe_dst_is_int_q[i] : mid_pipe_dst_is_int_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:389:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:389:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:389:187
					mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:389:295
					mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= (reg_ena ? mid_pipe_info_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 8+:8] : mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:390:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:390:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:390:187
					mid_pipe_mant_zero_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:390:295
					mid_pipe_mant_zero_q[i + 1] <= (reg_ena ? mid_pipe_mant_zero_q[i] : mid_pipe_mant_zero_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:391:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:391:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:391:187
					mid_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:391:295
					mid_pipe_op_mod_q[i + 1] <= (reg_ena ? mid_pipe_op_mod_q[i] : mid_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:392:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:392:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:392:199
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:392:307
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:393:99
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:393:155
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:393:211
					mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:393:319
					mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:394:99
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:394:155
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:394:211
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:394:319
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:395:100
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:395:156
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:395:212
					mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_87CC5(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:395:320
					mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= (reg_ena ? mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] : mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:396:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:396:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:396:197
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:396:305
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:397:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:397:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:397:187
					mid_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:397:295
					mid_pipe_mask_q[i + 1] <= (reg_ena ? mid_pipe_mask_q[i] : mid_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:398:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:398:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:398:197
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:398:305
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:401:3
	assign input_sign_q = mid_pipe_input_sign_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:402:3
	assign input_exp_q = mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:403:3
	assign input_mant_q = mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:404:3
	assign destination_exp_q = mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:405:3
	assign src_is_int_q = mid_pipe_src_is_int_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:406:3
	assign dst_is_int_q = mid_pipe_dst_is_int_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:407:3
	assign info_q = mid_pipe_info_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 8+:8];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:408:3
	assign mant_is_zero_q = mid_pipe_mant_zero_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:409:3
	assign op_mod_q2 = mid_pipe_op_mod_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:410:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:411:3
	assign src_fmt_q2 = mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:412:3
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:413:3
	assign int_fmt_q2 = mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:418:3
	reg [INT_EXP_WIDTH - 1:0] final_exp;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:420:3
	reg [2 * INT_MAN_WIDTH:0] preshift_mant;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:421:3
	wire [2 * INT_MAN_WIDTH:0] destination_mant;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:422:3
	wire [SUPER_MAN_BITS - 1:0] final_mant;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:423:3
	wire [MAX_INT_WIDTH - 1:0] final_int;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:425:3
	reg [$clog2(INT_MAN_WIDTH + 1) - 1:0] denorm_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:427:3
	wire [1:0] fp_round_sticky_bits;
	wire [1:0] int_round_sticky_bits;
	wire [1:0] round_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:428:3
	reg of_before_round;
	reg uf_before_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:432:3
	always @(*) begin : cast_value
		// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:434:5
		final_exp = $unsigned(destination_exp_q);
		// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:435:5
		preshift_mant = 1'sb0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:436:5
		denorm_shamt = SUPER_MAN_BITS - fpnew_pkg_man_bits(dst_fmt_q2);
		// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:437:5
		of_before_round = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:438:5
		uf_before_round = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:441:5
		preshift_mant = input_mant_q << (INT_MAN_WIDTH + 1);
		// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:444:5
		if (dst_is_int_q) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:446:7
			denorm_shamt = $unsigned((MAX_INT_WIDTH - 1) - input_exp_q);
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:448:7
			if ((input_exp_q >= $signed((fpnew_pkg_int_width(int_fmt_q2) - 1) + op_mod_q2)) && !(((!op_mod_q2 && input_sign_q) && (input_exp_q == $signed(fpnew_pkg_int_width(int_fmt_q2) - 1))) && (input_mant_q == {1'b1, {INT_MAN_WIDTH - 1 {1'b0}}}))) begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:453:9
				denorm_shamt = 1'sb0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:454:9
				of_before_round = 1'b1;
			end
			else if (input_exp_q < -1) begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:457:9
				denorm_shamt = MAX_INT_WIDTH + 1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:458:9
				uf_before_round = 1'b1;
			end
		end
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:463:7
			if ((destination_exp_q >= ($signed(2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1)) || (~src_is_int_q && info_q[4])) begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:465:9
				final_exp = $unsigned((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 2);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:466:9
				preshift_mant = 1'sb1;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:467:9
				of_before_round = 1'b1;
			end
			else if ((destination_exp_q < 1) && (destination_exp_q >= -$signed(fpnew_pkg_man_bits(dst_fmt_q2)))) begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:471:9
				final_exp = 1'sb0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:472:9
				denorm_shamt = $unsigned((denorm_shamt + 1) - destination_exp_q);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:473:9
				uf_before_round = 1'b1;
			end
			else if (destination_exp_q < -$signed(fpnew_pkg_man_bits(dst_fmt_q2))) begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:476:9
				final_exp = 1'sb0;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:477:9
				denorm_shamt = $unsigned((denorm_shamt + 2) + fpnew_pkg_man_bits(dst_fmt_q2));
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:478:9
				uf_before_round = 1'b1;
			end
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:483:3
	localparam NUM_FP_STICKY = ((2 * INT_MAN_WIDTH) - SUPER_MAN_BITS) - 1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:484:3
	localparam NUM_INT_STICKY = (2 * INT_MAN_WIDTH) - MAX_INT_WIDTH;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:487:3
	assign destination_mant = preshift_mant >> denorm_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:489:3
	assign {final_mant, fp_round_sticky_bits[1]} = destination_mant[(2 * INT_MAN_WIDTH) - 1-:SUPER_MAN_BITS + 1];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:491:3
	assign {final_int, int_round_sticky_bits[1]} = destination_mant[2 * INT_MAN_WIDTH-:MAX_INT_WIDTH + 1];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:493:3
	assign fp_round_sticky_bits[0] = |{destination_mant[NUM_FP_STICKY - 1:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:494:3
	assign int_round_sticky_bits[0] = |{destination_mant[NUM_INT_STICKY - 1:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:497:3
	assign round_sticky_bits = (dst_is_int_q ? int_round_sticky_bits : fp_round_sticky_bits);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:502:3
	wire [WIDTH - 1:0] pre_round_abs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:503:3
	wire of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:504:3
	wire uf_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:506:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_pre_round_abs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:507:3
	reg [4:0] fmt_of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:508:3
	reg [4:0] fmt_uf_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:510:3
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_pre_round_abs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:511:3
	reg [3:0] ifmt_of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:513:3
	wire rounded_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:514:3
	wire [WIDTH - 1:0] rounded_abs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:515:3
	wire result_true_zero;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:517:3
	wire [WIDTH - 1:0] rounded_int_res;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:518:3
	wire rounded_int_res_zero;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:522:3
	genvar _gv_fmt_10;
	generate
		for (_gv_fmt_10 = 0; _gv_fmt_10 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_10 = _gv_fmt_10 + 1) begin : gen_res_assemble
			localparam fmt = _gv_fmt_10;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:524:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:525:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:528:7
				always @(*) begin : assemble_result
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:529:9
					fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = {final_exp[EXP_BITS - 1:0], final_mant[MAN_BITS - 1:0]};
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:532:7
				wire [WIDTH * 1:1] sv2v_tmp_C33E0;
				assign sv2v_tmp_C33E0 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = sv2v_tmp_C33E0;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:537:3
	genvar _gv_ifmt_4;
	generate
		for (_gv_ifmt_4 = 0; _gv_ifmt_4 < sv2v_cast_32_signed(NUM_INT_FORMATS); _gv_ifmt_4 = _gv_ifmt_4 + 1) begin : gen_int_res_sign_ext
			localparam ifmt = _gv_ifmt_4;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:539:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:542:7
				always @(*) begin : assemble_result
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:544:9
					ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = {WIDTH {final_int[INT_WIDTH - 1]}};
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:545:9
					ifmt_pre_round_abs[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = final_int[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:548:7
				wire [WIDTH * 1:1] sv2v_tmp_F6FA8;
				assign sv2v_tmp_F6FA8 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = sv2v_tmp_F6FA8;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:553:3
	assign pre_round_abs = (dst_is_int_q ? ifmt_pre_round_abs[int_fmt_q2 * WIDTH+:WIDTH] : fmt_pre_round_abs[dst_fmt_q2 * WIDTH+:WIDTH]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:555:3
	fpnew_rounding #(.AbsWidth(WIDTH)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(input_sign_q),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(1'b0),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_true_zero)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:568:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:571:3
	genvar _gv_fmt_11;
	generate
		for (_gv_fmt_11 = 0; _gv_fmt_11 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_11 = _gv_fmt_11 + 1) begin : gen_sign_inject
			localparam fmt = _gv_fmt_11;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:573:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:574:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:575:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:578:7
				always @(*) begin : post_process
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:580:9
					fmt_uf_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:581:9
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:584:9
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:585:9
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = (src_is_int_q & mant_is_zero_q ? {FP_WIDTH * 1 {1'sb0}} : {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]});
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:590:7
				wire [1:1] sv2v_tmp_4A747;
				assign sv2v_tmp_4A747 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4A747;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:591:7
				wire [1:1] sv2v_tmp_90681;
				assign sv2v_tmp_90681 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_90681;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:592:7
				wire [WIDTH * 1:1] sv2v_tmp_649FB;
				assign sv2v_tmp_649FB = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_649FB;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:597:3
	assign rounded_int_res = (rounded_sign ? $unsigned(-rounded_abs) : rounded_abs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:598:3
	assign rounded_int_res_zero = rounded_int_res == {WIDTH {1'sb0}};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:601:3
	genvar _gv_ifmt_5;
	generate
		for (_gv_ifmt_5 = 0; _gv_ifmt_5 < sv2v_cast_32_signed(NUM_INT_FORMATS); _gv_ifmt_5 = _gv_ifmt_5 + 1) begin : gen_int_overflow
			localparam ifmt = _gv_ifmt_5;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:603:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:606:7
				always @(*) begin : detect_overflow
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:607:9
					ifmt_of_after_round[ifmt] = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:609:9
					if (!rounded_sign && (input_exp_q == $signed((INT_WIDTH - 2) + op_mod_q2)))
						// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:611:11
						ifmt_of_after_round[ifmt] = ~rounded_int_res[(INT_WIDTH - 2) + op_mod_q2];
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:615:7
				wire [1:1] sv2v_tmp_3841B;
				assign sv2v_tmp_3841B = fpnew_pkg_DONT_CARE;
				always @(*) ifmt_of_after_round[ifmt] = sv2v_tmp_3841B;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:620:3
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:621:3
	assign of_after_round = (dst_is_int_q ? ifmt_of_after_round[int_fmt_q2] : fmt_of_after_round[dst_fmt_q2]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:626:3
	wire [WIDTH - 1:0] fp_special_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:627:3
	wire [4:0] fp_special_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:628:3
	wire fp_result_is_special;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:630:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:633:3
	genvar _gv_fmt_12;
	generate
		for (_gv_fmt_12 = 0; _gv_fmt_12 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_12 = _gv_fmt_12 + 1) begin : gen_special_results
			localparam fmt = _gv_fmt_12;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:635:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:636:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:637:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:639:5
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:640:5
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:643:7
				always @(*) begin : special_results
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:644:9
					reg [FP_WIDTH - 1:0] special_res;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:645:9
					special_res = (info_q[5] ? input_sign_q << (FP_WIDTH - 1) : {1'b0, QNAN_EXPONENT, QNAN_MANTISSA});
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:650:9
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:651:9
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:654:7
				wire [WIDTH * 1:1] sv2v_tmp_B718F;
				assign sv2v_tmp_B718F = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_B718F;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:659:3
	assign fp_result_is_special = ~src_is_int_q & ((info_q[5] | info_q[3]) | ~info_q[0]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:664:3
	assign fp_special_status = {info_q[2], 4'b0000};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:667:3
	assign fp_special_result = fmt_special_result[dst_fmt_q2 * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:672:3
	wire [WIDTH - 1:0] int_special_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:673:3
	wire [4:0] int_special_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:674:3
	wire int_result_is_special;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:676:3
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_special_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:679:3
	genvar _gv_ifmt_6;
	generate
		for (_gv_ifmt_6 = 0; _gv_ifmt_6 < sv2v_cast_32_signed(NUM_INT_FORMATS); _gv_ifmt_6 = _gv_ifmt_6 + 1) begin : gen_special_results_int
			localparam ifmt = _gv_ifmt_6;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:681:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:684:7
				always @(*) begin : special_results
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:685:9
					reg [INT_WIDTH - 1:0] special_res;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:688:9
					special_res[INT_WIDTH - 2:0] = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:689:9
					special_res[INT_WIDTH - 1] = op_mod_q2;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:692:9
					if (input_sign_q && !info_q[3])
						// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:693:11
						special_res = ~special_res;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:696:9
					ifmt_special_result[ifmt * WIDTH+:WIDTH] = {WIDTH {special_res[INT_WIDTH - 1]}};
					// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:697:9
					ifmt_special_result[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:700:7
				wire [WIDTH * 1:1] sv2v_tmp_99B6D;
				assign sv2v_tmp_99B6D = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_special_result[ifmt * WIDTH+:WIDTH] = sv2v_tmp_99B6D;
			end
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:705:3
	assign int_result_is_special = ((((info_q[3] | info_q[4]) | of_before_round) | of_after_round) | ~info_q[0]) | ((input_sign_q & op_mod_q2) & ~rounded_int_res_zero);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:710:3
	assign int_special_status = 5'b10000;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:713:3
	assign int_special_result = ifmt_special_result[int_fmt_q2 * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:718:3
	wire [4:0] int_regular_status;
	wire [4:0] fp_regular_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:720:3
	wire [WIDTH - 1:0] fp_result;
	wire [WIDTH - 1:0] int_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:721:3
	wire [4:0] fp_status;
	wire [4:0] int_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:723:3
	assign fp_regular_status[4] = src_is_int_q & (of_before_round | of_after_round);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:724:3
	assign fp_regular_status[3] = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:725:3
	assign fp_regular_status[2] = ~src_is_int_q & (~info_q[4] & (of_before_round | of_after_round));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:726:3
	assign fp_regular_status[1] = uf_after_round & fp_regular_status[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:727:3
	assign fp_regular_status[0] = (src_is_int_q ? |fp_round_sticky_bits : |fp_round_sticky_bits | (~info_q[4] & (of_before_round | of_after_round)));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:729:3
	assign int_regular_status = {4'b0000, |int_round_sticky_bits};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:731:3
	assign fp_result = (fp_result_is_special ? fp_special_result : fmt_result[dst_fmt_q2 * WIDTH+:WIDTH]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:732:3
	assign fp_status = (fp_result_is_special ? fp_special_status : fp_regular_status);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:733:3
	assign int_result = (int_result_is_special ? int_special_result : rounded_int_res);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:734:3
	assign int_status = (int_result_is_special ? int_special_status : int_regular_status);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:737:3
	wire [WIDTH - 1:0] result_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:738:3
	wire [4:0] status_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:739:3
	wire extension_bit;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:742:3
	assign result_d = (dst_is_int_q ? int_result : fp_result);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:743:3
	assign status_d = (dst_is_int_q ? int_status : fp_status);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:746:3
	assign extension_bit = (dst_is_int_q ? int_result[WIDTH - 1] : 1'b1);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:752:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:753:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:754:3
	reg [0:NUM_OUT_REGS] out_pipe_ext_bit_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:755:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] out_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:756:3
	reg [0:NUM_OUT_REGS] out_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:757:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:758:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:760:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:763:3
	wire [WIDTH * 1:1] sv2v_tmp_4086F;
	assign sv2v_tmp_4086F = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_4086F;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:764:3
	wire [5:1] sv2v_tmp_B7C45;
	assign sv2v_tmp_B7C45 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_B7C45;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:765:3
	wire [1:1] sv2v_tmp_8F736;
	assign sv2v_tmp_8F736 = extension_bit;
	always @(*) out_pipe_ext_bit_q[0] = sv2v_tmp_8F736;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:766:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_A76BD;
	assign sv2v_tmp_A76BD = mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_A76BD;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:767:3
	wire [1:1] sv2v_tmp_DB780;
	assign sv2v_tmp_DB780 = mid_pipe_mask_q[NUM_MID_REGS];
	always @(*) out_pipe_mask_q[0] = sv2v_tmp_DB780;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:768:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_17955;
	assign sv2v_tmp_17955 = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_17955;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:769:3
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:771:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:773:3
	genvar _gv_i_230;
	generate
		for (_gv_i_230 = 0; _gv_i_230 < NUM_OUT_REGS; _gv_i_230 = _gv_i_230 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_230;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:775:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:779:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:781:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:781:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:781:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:781:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:783:5
			assign reg_ena = (out_pipe_ready[i] & out_pipe_valid_q[i]) | reg_ena_i[(NUM_INP_REGS + NUM_MID_REGS) + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:785:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:785:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:785:181
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:785:289
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:786:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:786:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:786:181
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:786:289
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:787:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:787:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:787:181
					out_pipe_ext_bit_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:787:289
					out_pipe_ext_bit_q[i + 1] <= (reg_ena ? out_pipe_ext_bit_q[i] : out_pipe_ext_bit_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:788:79
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:788:135
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:788:191
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:788:299
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:789:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:789:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:789:181
					out_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:789:289
					out_pipe_mask_q[i + 1] <= (reg_ena ? out_pipe_mask_q[i] : out_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:790:79
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:790:135
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:790:191
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:790:299
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:793:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:795:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:796:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:797:3
	assign extension_bit_o = out_pipe_ext_bit_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:798:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:799:3
	assign mask_o = out_pipe_mask_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:800:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:801:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_cast_multi.sv:802:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_noncomp_59FAB_0570D (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	mask_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	class_mask_o,
	is_class_o,
	tag_o,
	mask_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o,
	reg_ena_i
);
	// removed localparam type TagType_TagType_TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:19:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:20:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:21:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:22:38
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:23:38
	// removed localparam type AuxType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:25:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:26:14
	localparam [31:0] ExtRegEnaWidth = (NumPipeRegs == 0 ? 1 : NumPipeRegs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:28:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:29:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:31:3
	input wire [(2 * WIDTH) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:32:3
	input wire [1:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:33:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:34:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:35:3
	input wire op_mod_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:36:3
	input wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:37:3
	input wire mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:38:3
	input wire aux_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:40:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:41:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:42:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:44:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:45:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:46:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:47:3
	// removed localparam type fpnew_pkg_classmask_e
	output wire [9:0] class_mask_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:48:3
	output wire is_class_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:49:3
	output wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:50:3
	output wire mask_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:51:3
	output wire aux_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:53:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:54:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:56:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:58:3
	input wire [ExtRegEnaWidth - 1:0] reg_ena_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:64:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:337:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:338:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:65:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:342:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:343:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:67:3
	localparam NUM_INP_REGS = ((PipeConfig == 2'd0) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:72:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:81:3
	// removed localparam type fp_t
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:91:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:92:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)] inp_pipe_is_boxed_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:93:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:94:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:95:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:96:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] inp_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:97:3
	reg [0:NUM_INP_REGS] inp_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:98:3
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:99:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:101:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:104:3
	wire [2 * WIDTH:1] sv2v_tmp_D1067;
	assign sv2v_tmp_D1067 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_D1067;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:105:3
	wire [2:1] sv2v_tmp_86D63;
	assign sv2v_tmp_86D63 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2+:2] = sv2v_tmp_86D63;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:106:3
	wire [3:1] sv2v_tmp_62109;
	assign sv2v_tmp_62109 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_62109;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:107:3
	wire [4:1] sv2v_tmp_0B797;
	assign sv2v_tmp_0B797 = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_0B797;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:108:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:109:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_622E2;
	assign sv2v_tmp_622E2 = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_622E2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:110:3
	wire [1:1] sv2v_tmp_407DF;
	assign sv2v_tmp_407DF = mask_i;
	always @(*) inp_pipe_mask_q[0] = sv2v_tmp_407DF;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:111:3
	wire [1:1] sv2v_tmp_8D189;
	assign sv2v_tmp_8D189 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_8D189;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:112:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:114:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:116:3
	genvar _gv_i_231;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] sv2v_cast_48BE4;
		input reg [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] inp;
		sv2v_cast_48BE4 = inp;
	endfunction
	generate
		for (_gv_i_231 = 0; _gv_i_231 < NUM_INP_REGS; _gv_i_231 = _gv_i_231 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_231;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:118:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:122:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:124:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:124:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:124:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:124:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:126:5
			assign reg_ena = (inp_pipe_ready[i] & inp_pipe_valid_q[i]) | reg_ena_i[i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:128:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:128:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:128:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:128:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:129:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:129:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:129:183
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:129:291
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2+:2] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:130:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:130:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:130:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:130:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:131:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:131:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:131:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:131:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:132:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:132:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:132:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:132:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:133:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:133:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:133:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:133:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:134:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:134:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:134:183
					inp_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:134:291
					inp_pipe_mask_q[i + 1] <= (reg_ena ? inp_pipe_mask_q[i] : inp_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:135:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:135:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:135:193
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:135:301
					inp_pipe_aux_q[i + 1] <= (reg_ena ? inp_pipe_aux_q[i] : inp_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:141:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [15:0] info_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:144:3
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(2)
	) i_class_a(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2+:2]),
		.info_o(info_q)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:153:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:154:3
	wire [7:0] info_a;
	wire [7:0] info_b;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:157:3
	assign operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:158:3
	assign operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:159:3
	assign info_a = info_q[0+:8];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:160:3
	assign info_b = info_q[8+:8];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:162:3
	wire any_operand_inf;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:163:3
	wire any_operand_nan;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:164:3
	wire signalling_nan;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:167:3
	assign any_operand_inf = |{info_a[4], info_b[4]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:168:3
	assign any_operand_nan = |{info_a[3], info_b[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:169:3
	assign signalling_nan = |{info_a[2], info_b[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:171:3
	wire operands_equal;
	wire operand_a_smaller;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:174:3
	assign operands_equal = (operand_a == operand_b) || (info_a[5] && info_b[5]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:176:3
	assign operand_a_smaller = (operand_a < operand_b) ^ (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] || operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:181:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] sgnj_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:182:3
	wire [4:0] sgnj_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:183:3
	wire sgnj_extension_bit;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:187:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_F2D56;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_F2D56 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_14681;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_14681 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_91364;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_91364 = inp;
	endfunction
	always @(*) begin : sign_injections
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:188:5
		reg sign_a;
		reg sign_b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:190:5
		sgnj_result = operand_a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:193:5
		if (!info_a[0])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:193:27
			sgnj_result = {1'b0, sv2v_cast_F2D56(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:196:5
		sign_a = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] & info_a[0];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:197:5
		sign_b = operand_b[1 + (EXP_BITS + (MAN_BITS - 1))] & info_b[0];
		case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
			3'b000:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:201:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_b;
			3'b001:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:202:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = ~sign_b;
			3'b010:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:203:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_a ^ sign_b;
			3'b011:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:204:23
				sgnj_result = operand_a;
			default:
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:205:16
				sgnj_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
		endcase
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:209:3
	assign sgnj_status = 1'sb0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:212:3
	assign sgnj_extension_bit = (inp_pipe_op_mod_q[NUM_INP_REGS] ? sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] : 1'b1);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:217:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] minmax_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:218:3
	reg [4:0] minmax_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:219:3
	wire minmax_extension_bit;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:223:3
	always @(*) begin : min_max
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:225:5
		minmax_status = 1'sb0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:228:5
		minmax_status[4] = signalling_nan;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:231:5
		if (info_a[3] && info_b[3])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:232:7
			minmax_result = {1'b0, sv2v_cast_F2D56(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		else if (info_a[3])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:234:29
			minmax_result = operand_b;
		else if (info_b[3])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:235:29
			minmax_result = operand_a;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:238:7
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000:
					// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:239:25
					minmax_result = (operand_a_smaller ? operand_a : operand_b);
				3'b001:
					// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:240:25
					minmax_result = (operand_a_smaller ? operand_b : operand_a);
				default:
					// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:241:18
					minmax_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
			endcase
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:246:3
	assign minmax_extension_bit = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:251:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] cmp_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:252:3
	reg [4:0] cmp_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:253:3
	wire cmp_extension_bit;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:258:3
	always @(*) begin : comparisons
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:260:5
		cmp_result = 1'sb0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:261:5
		cmp_status = 1'sb0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:264:5
		if (signalling_nan) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:265:7
			cmp_status[4] = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:266:7
			cmp_result = (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3] == 3'b010) && inp_pipe_op_mod_q[NUM_INP_REGS];
		end
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:269:7
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000:
					// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:271:11
					if (any_operand_nan)
						// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:271:32
						cmp_status[4] = 1'b1;
					else
						// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:272:16
						cmp_result = (operand_a_smaller | operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b001:
					// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:275:11
					if (any_operand_nan)
						// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:275:32
						cmp_status[4] = 1'b1;
					else
						// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:276:16
						cmp_result = (operand_a_smaller & ~operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b010:
					// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:279:11
					if (any_operand_nan)
						// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:279:32
						cmp_result = inp_pipe_op_mod_q[NUM_INP_REGS];
					else
						// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:280:16
						cmp_result = operands_equal ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				default:
					// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:282:18
					cmp_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
			endcase
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:287:3
	assign cmp_extension_bit = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:292:3
	wire [4:0] class_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:293:3
	wire class_extension_bit;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:294:3
	reg [9:0] class_mask_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:297:3
	always @(*) begin : classify
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:298:5
		if (info_a[7])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:299:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000010 : 10'b0001000000);
		else if (info_a[6])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:301:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000100 : 10'b0000100000);
		else if (info_a[5])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:303:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000001000 : 10'b0000010000);
		else if (info_a[4])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:305:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000001 : 10'b0010000000);
		else if (info_a[3])
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:307:7
			class_mask_d = (info_a[2] ? 10'b0100000000 : 10'b1000000000);
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:309:7
			class_mask_d = 10'b1000000000;
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:313:3
	assign class_status = 1'sb0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:314:3
	assign class_extension_bit = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:319:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:320:3
	reg [4:0] status_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:321:3
	reg extension_bit_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:322:3
	wire is_class_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:325:3
	always @(*) begin : select_result
		// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:326:5
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(6): begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:328:9
				result_d = sgnj_result;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:329:9
				status_d = sgnj_status;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:330:9
				extension_bit_d = sgnj_extension_bit;
			end
			sv2v_cast_A53F3(7): begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:333:9
				result_d = minmax_result;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:334:9
				status_d = minmax_status;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:335:9
				extension_bit_d = minmax_extension_bit;
			end
			sv2v_cast_A53F3(8): begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:338:9
				result_d = cmp_result;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:339:9
				status_d = cmp_status;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:340:9
				extension_bit_d = cmp_extension_bit;
			end
			sv2v_cast_A53F3(9): begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:343:9
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:344:9
				status_d = class_status;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:345:9
				extension_bit_d = class_extension_bit;
			end
			default: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:348:9
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:349:9
				status_d = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:350:9
				extension_bit_d = fpnew_pkg_DONT_CARE;
			end
		endcase
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:355:3
	assign is_class_d = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(9);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:361:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:362:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:363:3
	reg [0:NUM_OUT_REGS] out_pipe_extension_bit_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:364:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 10) + ((NUM_OUT_REGS * 10) - 1) : ((NUM_OUT_REGS + 1) * 10) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 10 : 0)] out_pipe_class_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:365:3
	reg [0:NUM_OUT_REGS] out_pipe_is_class_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:366:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] out_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:367:3
	reg [0:NUM_OUT_REGS] out_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:368:3
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:369:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:371:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:374:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_07494;
	assign sv2v_tmp_07494 = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_07494;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:375:3
	wire [5:1] sv2v_tmp_CCE43;
	assign sv2v_tmp_CCE43 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_CCE43;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:376:3
	wire [1:1] sv2v_tmp_8E9A9;
	assign sv2v_tmp_8E9A9 = extension_bit_d;
	always @(*) out_pipe_extension_bit_q[0] = sv2v_tmp_8E9A9;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:377:3
	wire [10:1] sv2v_tmp_94259;
	assign sv2v_tmp_94259 = class_mask_d;
	always @(*) out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 10+:10] = sv2v_tmp_94259;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:378:3
	wire [1:1] sv2v_tmp_7DF01;
	assign sv2v_tmp_7DF01 = is_class_d;
	always @(*) out_pipe_is_class_q[0] = sv2v_tmp_7DF01;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:379:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_0F5B6;
	assign sv2v_tmp_0F5B6 = inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_0F5B6;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:380:3
	wire [1:1] sv2v_tmp_20A3C;
	assign sv2v_tmp_20A3C = inp_pipe_mask_q[NUM_INP_REGS];
	always @(*) out_pipe_mask_q[0] = sv2v_tmp_20A3C;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:381:3
	wire [1:1] sv2v_tmp_FA930;
	assign sv2v_tmp_FA930 = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_FA930;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:382:3
	wire [1:1] sv2v_tmp_2CB8C;
	assign sv2v_tmp_2CB8C = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_2CB8C;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:384:3
	assign inp_pipe_ready[NUM_INP_REGS] = out_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:386:3
	genvar _gv_i_232;
	generate
		for (_gv_i_232 = 0; _gv_i_232 < NUM_OUT_REGS; _gv_i_232 = _gv_i_232 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_232;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:388:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:392:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:394:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:394:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:394:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:394:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:396:5
			assign reg_ena = (out_pipe_ready[i] & out_pipe_valid_q[i]) | reg_ena_i[NUM_INP_REGS + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:398:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:398:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:398:193
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:398:301
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:399:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:399:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:399:193
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:399:301
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:400:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:400:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:400:193
					out_pipe_extension_bit_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:400:301
					out_pipe_extension_bit_q[i + 1] <= (reg_ena ? out_pipe_extension_bit_q[i] : out_pipe_extension_bit_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:401:94
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:401:150
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:401:206
					out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= 10'b1000000000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:401:314
					out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= (reg_ena ? out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 10+:10] : out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:402:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:402:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:402:193
					out_pipe_is_class_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:402:301
					out_pipe_is_class_q[i + 1] <= (reg_ena ? out_pipe_is_class_q[i] : out_pipe_is_class_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:403:91
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:403:147
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:403:203
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:403:311
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:404:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:404:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:404:193
					out_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:404:301
					out_pipe_mask_q[i + 1] <= (reg_ena ? out_pipe_mask_q[i] : out_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:405:91
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:405:147
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:405:203
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:405:311
					out_pipe_aux_q[i + 1] <= (reg_ena ? out_pipe_aux_q[i] : out_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:408:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:410:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:411:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:412:3
	assign extension_bit_o = out_pipe_extension_bit_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:413:3
	assign class_mask_o = out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 10+:10];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:414:3
	assign is_class_o = out_pipe_is_class_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:415:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:416:3
	assign mask_o = out_pipe_mask_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:417:3
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:418:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_noncomp.sv:419:3
	assign busy_o = |{inp_pipe_valid_q, out_pipe_valid_q};
endmodule
// removed package "fpnew_pkg"
module fpnew_classifier (
	operands_i,
	is_boxed_i,
	info_o
);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:18:13
	parameter [31:0] NumOperands = 1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:20:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:22:3
	input wire [(NumOperands * WIDTH) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:23:3
	input wire [NumOperands - 1:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:24:3
	// removed localparam type fpnew_pkg_fp_info_t
	output reg [(NumOperands * 8) - 1:0] info_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:27:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:337:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:338:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:28:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:342:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:343:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:31:3
	// removed localparam type fp_t
	// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:38:3
	genvar _gv_op_3;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_op_3 = 0; _gv_op_3 < sv2v_cast_32_signed(NumOperands); _gv_op_3 = _gv_op_3 + 1) begin : gen_num_values
			localparam op = _gv_op_3;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:40:5
			reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] value;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:41:5
			reg is_boxed;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:42:5
			reg is_normal;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:43:5
			reg is_inf;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:44:5
			reg is_nan;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:45:5
			reg is_signalling;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:46:5
			reg is_quiet;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:47:5
			reg is_zero;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:48:5
			reg is_subnormal;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:53:5
			always @(*) begin : classify_input
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:54:7
				value = operands_i[op * WIDTH+:WIDTH];
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:55:7
				is_boxed = is_boxed_i[op];
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:56:7
				is_normal = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] != {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] != {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}});
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:57:7
				is_zero = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && (value[MAN_BITS - 1-:MAN_BITS] == {MAN_BITS * 1 {1'sb0}});
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:58:7
				is_subnormal = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && !is_zero;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:59:7
				is_inf = is_boxed && ((value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}}) && (value[MAN_BITS - 1-:MAN_BITS] == {MAN_BITS * 1 {1'sb0}}));
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:60:7
				is_nan = !is_boxed || ((value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}}) && (value[MAN_BITS - 1-:MAN_BITS] != {MAN_BITS * 1 {1'sb0}}));
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:61:7
				is_signalling = (is_boxed && is_nan) && (value[(MAN_BITS - 1) - ((MAN_BITS - 1) - (MAN_BITS - 1))] == 1'b0);
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:62:7
				is_quiet = is_nan && !is_signalling;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:64:7
				info_o[(op * 8) + 7] = is_normal;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:65:7
				info_o[(op * 8) + 6] = is_subnormal;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:66:7
				info_o[(op * 8) + 5] = is_zero;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:67:7
				info_o[(op * 8) + 4] = is_inf;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:68:7
				info_o[(op * 8) + 3] = is_nan;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:69:7
				info_o[(op * 8) + 2] = is_signalling;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:70:7
				info_o[(op * 8) + 1] = is_quiet;
				// Trace: /vortex/third_party/cvfpu/src/fpnew_classifier.sv:71:7
				info_o[op * 8] = is_boxed;
			end
		end
	endgenerate
endmodule
module fpnew_fma_7C8F3_7759B (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	mask_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	mask_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o,
	reg_ena_i
);
	// removed localparam type TagType_TagType_TagType_TagType_TAG_WIDTH_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAG_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:19:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:20:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:21:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:22:38
	// removed localparam type TagType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:23:38
	// removed localparam type AuxType
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:25:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:314:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:315:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:26:14
	localparam [31:0] ExtRegEnaWidth = (NumPipeRegs == 0 ? 1 : NumPipeRegs);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:28:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:29:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:31:3
	input wire [(3 * WIDTH) - 1:0] operands_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:32:3
	input wire [2:0] is_boxed_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:33:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:34:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:35:3
	input wire op_mod_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:36:3
	input wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:37:3
	input wire mask_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:38:3
	input wire aux_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:40:3
	input wire in_valid_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:41:3
	output wire in_ready_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:42:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:44:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:45:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:46:3
	output wire extension_bit_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:47:3
	output wire [TagType_TagType_TagType_TagType_TAG_WIDTH + 0:0] tag_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:48:3
	output wire mask_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:49:3
	output wire aux_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:51:3
	output wire out_valid_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:52:3
	input wire out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:54:3
	output wire busy_o;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:56:3
	input wire [ExtRegEnaWidth - 1:0] reg_ena_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:62:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:337:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:338:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:63:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:342:44
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:343:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:64:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:347:40
		input reg [2:0] fmt;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:348:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	localparam [31:0] BIAS = fpnew_pkg_bias(FpFormat);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:66:3
	localparam [31:0] PRECISION_BITS = MAN_BITS + 1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:68:3
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:69:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:73:3
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:34
		input reg signed [31:0] a;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:306:41
		input reg signed [31:0] b;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_pkg.sv:307:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	localparam [31:0] EXP_WIDTH = $unsigned(fpnew_pkg_maximum(EXP_BITS + 2, LZC_RESULT_WIDTH));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:75:3
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 5);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:77:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:82:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:87:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:96:3
	// removed localparam type fp_t
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:106:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:107:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_is_boxed_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:108:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:109:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:110:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:111:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] inp_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:112:3
	reg [0:NUM_INP_REGS] inp_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:113:3
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:114:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:116:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:119:3
	wire [3 * WIDTH:1] sv2v_tmp_BC8B9;
	assign sv2v_tmp_BC8B9 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_BC8B9;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:120:3
	wire [3:1] sv2v_tmp_FE389;
	assign sv2v_tmp_FE389 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_FE389;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:121:3
	wire [3:1] sv2v_tmp_E1339;
	assign sv2v_tmp_E1339 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_E1339;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:122:3
	wire [4:1] sv2v_tmp_CBA8F;
	assign sv2v_tmp_CBA8F = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_CBA8F;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:123:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:124:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_FAE22;
	assign sv2v_tmp_FAE22 = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_FAE22;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:125:3
	wire [1:1] sv2v_tmp_407DF;
	assign sv2v_tmp_407DF = mask_i;
	always @(*) inp_pipe_mask_q[0] = sv2v_tmp_407DF;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:126:3
	wire [1:1] sv2v_tmp_8D189;
	assign sv2v_tmp_8D189 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_8D189;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:127:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:129:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:131:3
	genvar _gv_i_233;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] sv2v_cast_48BE4;
		input reg [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) - 1:0] inp;
		sv2v_cast_48BE4 = inp;
	endfunction
	generate
		for (_gv_i_233 = 0; _gv_i_233 < NUM_INP_REGS; _gv_i_233 = _gv_i_233 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_233;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:133:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:137:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:139:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:139:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:139:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:139:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:141:5
			assign reg_ena = (inp_pipe_ready[i] & inp_pipe_valid_q[i]) | reg_ena_i[i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:143:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:143:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:143:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:143:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:144:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:144:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:144:183
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:144:291
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:145:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:145:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:145:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:145:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:146:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:146:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:146:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:146:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:147:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:147:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:147:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:147:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:148:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:148:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:148:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:148:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:149:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:149:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:149:183
					inp_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:149:291
					inp_pipe_mask_q[i + 1] <= (reg_ena ? inp_pipe_mask_q[i] : inp_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:150:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:150:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:150:193
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:150:301
					inp_pipe_aux_q[i + 1] <= (reg_ena ? inp_pipe_aux_q[i] : inp_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:156:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [23:0] info_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:159:3
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(3)
	) i_class_inputs(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3]),
		.info_o(info_q)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:168:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_c;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:169:3
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:183:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_91364;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_91364 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_60B87;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_60B87 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_F33EE;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_F33EE = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_14681;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_14681 = inp;
	endfunction
	always @(*) begin : op_select
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:186:5
		operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:187:5
		operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:188:5
		operand_c = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:189:5
		info_a = info_q[0+:8];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:190:5
		info_b = info_q[8+:8];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:191:5
		info_c = info_q[16+:8];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:194:5
		operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] = operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:196:5
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(0):
				;
			sv2v_cast_A53F3(1):
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:198:26
				operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] = ~operand_a[1 + (EXP_BITS + (MAN_BITS - 1))];
			sv2v_cast_A53F3(2), sv2v_cast_A53F3(15): begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:201:9
				operand_a = {1'b0, sv2v_cast_91364(BIAS), sv2v_cast_60B87(1'sb0)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:202:9
				info_a = 8'b10000001;
			end
			sv2v_cast_A53F3(3): begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:205:9
				if (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3] == 3'b010)
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:206:11
					operand_c = {1'b0, sv2v_cast_F33EE(1'sb0), sv2v_cast_60B87(1'sb0)};
				else
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:208:11
					operand_c = {1'b1, sv2v_cast_F33EE(1'sb0), sv2v_cast_60B87(1'sb0)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:209:9
				info_c = 8'b00100001;
			end
			default: begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:212:9
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:213:9
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:214:9
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:215:9
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:216:9
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:217:9
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:225:3
	wire any_operand_inf;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:226:3
	wire any_operand_nan;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:227:3
	wire signalling_nan;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:228:3
	wire effective_subtraction;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:229:3
	wire tentative_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:232:3
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:233:3
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:234:3
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:236:3
	assign effective_subtraction = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]) ^ operand_c[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:238:3
	assign tentative_sign = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:243:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:244:3
	reg [4:0] special_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:245:3
	reg result_is_special;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:247:3
	always @(*) begin : special_cases
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:249:5
		special_result = {1'b0, sv2v_cast_F33EE(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:250:5
		special_status = 1'sb0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:251:5
		result_is_special = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:257:5
		if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:258:7
			result_is_special = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:259:7
			special_status[4] = 1'b1;
		end
		else if (any_operand_nan) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:262:7
			result_is_special = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:263:7
			special_status[4] = signalling_nan;
		end
		else if (any_operand_inf) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:266:7
			result_is_special = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:268:7
			if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:269:9
				special_status[4] = 1'b1;
			else if (info_a[4] || info_b[4])
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:273:9
				special_result = {operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_F33EE(1'sb1), sv2v_cast_60B87(1'sb0)};
			else if (info_c[4])
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:277:9
				special_result = {operand_c[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_F33EE(1'sb1), sv2v_cast_60B87(1'sb0)};
		end
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:285:3
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:286:3
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:287:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:290:3
	assign exponent_a = $signed({1'b0, operand_a[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:291:3
	assign exponent_b = $signed({1'b0, operand_b[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:292:3
	assign exponent_c = $signed({1'b0, operand_c[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:296:3
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:298:3
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(BIAS) : $signed((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - $signed(BIAS)));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:304:3
	assign exponent_difference = exponent_addend - exponent_product;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:306:3
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:309:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:311:3
	always @(*) begin : addend_shift_amount
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:313:5
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:314:7
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:317:7
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:320:7
			addend_shamt = 0;
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:326:3
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:327:3
	wire [(2 * PRECISION_BITS) - 1:0] product;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:328:3
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:331:3
	assign mantissa_a = {info_a[7], operand_a[MAN_BITS - 1-:MAN_BITS]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:332:3
	assign mantissa_b = {info_b[7], operand_b[MAN_BITS - 1-:MAN_BITS]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:333:3
	assign mantissa_c = {info_c[7], operand_c[MAN_BITS - 1-:MAN_BITS]};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:336:3
	assign product = mantissa_a * mantissa_b;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:341:3
	assign product_shifted = product << 2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:346:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:347:3
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:348:3
	wire sticky_before_add;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:349:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:350:3
	wire inject_carry_in;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:360:3
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:363:3
	assign sticky_before_add = |addend_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:367:3
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:368:3
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:373:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_pos;
	wire [(3 * PRECISION_BITS) + 4:0] sum_neg;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:374:3
	wire sum_carry;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:375:3
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:376:3
	wire final_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:379:3
	assign sum_pos = (product_shifted + addend_shifted) + inject_carry_in;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:380:3
	assign sum_carry = sum_pos[(3 * PRECISION_BITS) + 4];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:385:3
	assign sum_neg = addend_after_shift - product_shifted;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:388:3
	assign sum = (effective_subtraction && ~sum_carry ? sum_neg : sum_pos);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:391:3
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:399:3
	wire effective_subtraction_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:400:3
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:401:3
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:402:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:403:3
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:404:3
	wire sticky_before_add_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:405:3
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:406:3
	wire final_sign_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:407:3
	wire [2:0] rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:408:3
	wire result_is_special_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:409:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:410:3
	wire [4:0] special_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:412:3
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:413:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:414:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:415:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:416:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:417:3
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:418:3
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:419:3
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:420:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:421:3
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:422:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] mid_pipe_spec_res_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:423:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:424:3
	reg [(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_MID_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_MID_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_MID_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_MID_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] mid_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:425:3
	reg [0:NUM_MID_REGS] mid_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:426:3
	reg [0:NUM_MID_REGS] mid_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:427:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:429:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:432:3
	wire [1:1] sv2v_tmp_56A72;
	assign sv2v_tmp_56A72 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_56A72;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:433:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_2D21E;
	assign sv2v_tmp_2D21E = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_2D21E;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:434:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_00793;
	assign sv2v_tmp_00793 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_00793;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:435:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_B4C85;
	assign sv2v_tmp_B4C85 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_B4C85;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:436:3
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_83404;
	assign sv2v_tmp_83404 = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_83404;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:437:3
	wire [1:1] sv2v_tmp_6F5F7;
	assign sv2v_tmp_6F5F7 = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6F5F7;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:438:3
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_CEAB3;
	assign sv2v_tmp_CEAB3 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_CEAB3;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:439:3
	wire [1:1] sv2v_tmp_D7BD0;
	assign sv2v_tmp_D7BD0 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_D7BD0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:440:3
	wire [3:1] sv2v_tmp_A74E2;
	assign sv2v_tmp_A74E2 = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_A74E2;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:441:3
	wire [1:1] sv2v_tmp_7DEC5;
	assign sv2v_tmp_7DEC5 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_7DEC5;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:442:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_4A83E;
	assign sv2v_tmp_4A83E = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_4A83E;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:443:3
	wire [5:1] sv2v_tmp_EC01B;
	assign sv2v_tmp_EC01B = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_EC01B;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:444:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_AEEB4;
	assign sv2v_tmp_AEEB4 = inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	always @(*) mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_AEEB4;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:445:3
	wire [1:1] sv2v_tmp_D7646;
	assign sv2v_tmp_D7646 = inp_pipe_mask_q[NUM_INP_REGS];
	always @(*) mid_pipe_mask_q[0] = sv2v_tmp_D7646;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:446:3
	wire [1:1] sv2v_tmp_CDA0E;
	assign sv2v_tmp_CDA0E = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) mid_pipe_aux_q[0] = sv2v_tmp_CDA0E;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:447:3
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:449:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:452:3
	genvar _gv_i_234;
	generate
		for (_gv_i_234 = 0; _gv_i_234 < NUM_MID_REGS; _gv_i_234 = _gv_i_234 + 1) begin : gen_inside_pipeline
			localparam i = _gv_i_234;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:454:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:458:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:460:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:460:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:460:408
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:460:560
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:462:5
			assign reg_ena = (mid_pipe_ready[i] & mid_pipe_valid_q[i]) | reg_ena_i[NUM_INP_REGS + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:464:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:464:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:464:189
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:464:297
					mid_pipe_eff_sub_q[i + 1] <= (reg_ena ? mid_pipe_eff_sub_q[i] : mid_pipe_eff_sub_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:465:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:465:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:465:189
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:465:297
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:466:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:466:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:466:189
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:466:297
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:467:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:467:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:467:189
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:467:297
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:468:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:468:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:468:189
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:468:297
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= (reg_ena ? mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] : mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:469:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:469:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:469:189
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:469:297
					mid_pipe_sticky_q[i + 1] <= (reg_ena ? mid_pipe_sticky_q[i] : mid_pipe_sticky_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:470:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:470:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:470:189
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:470:297
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= (reg_ena ? mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] : mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:471:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:471:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:471:189
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:471:297
					mid_pipe_final_sign_q[i + 1] <= (reg_ena ? mid_pipe_final_sign_q[i] : mid_pipe_final_sign_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:472:89
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:472:145
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:472:201
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:472:309
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:473:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:473:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:473:189
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:473:297
					mid_pipe_res_is_spec_q[i + 1] <= (reg_ena ? mid_pipe_res_is_spec_q[i] : mid_pipe_res_is_spec_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:474:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:474:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:474:189
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:474:297
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:475:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:475:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:475:189
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:475:297
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= (reg_ena ? mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5] : mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:476:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:476:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:476:199
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:476:307
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:477:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:477:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:477:189
					mid_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:477:297
					mid_pipe_mask_q[i + 1] <= (reg_ena ? mid_pipe_mask_q[i] : mid_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:478:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:478:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:478:199
					mid_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:478:307
					mid_pipe_aux_q[i + 1] <= (reg_ena ? mid_pipe_aux_q[i] : mid_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:481:3
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:482:3
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:483:3
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:484:3
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:485:3
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:486:3
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:487:3
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:488:3
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:489:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:490:3
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:491:3
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:492:3
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:497:3
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:498:3
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:499:3
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:500:3
	wire lzc_zeroes;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:502:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:503:3
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:505:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:506:3
	reg [PRECISION_BITS:0] final_mantissa;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:507:3
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:508:3
	wire sticky_after_norm;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:510:3
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:512:3
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:515:3
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:524:3
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:527:3
	always @(*) begin : norm_shift_amount
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:529:5
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			begin
				// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:531:7
				if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:533:9
					norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:534:9
					normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
				end
				else begin
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:538:9
					norm_shamt = $unsigned(($signed(PRECISION_BITS) + 2) + exponent_product_q);
					// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:539:9
					normalized_exponent = 0;
				end
			end
		end
		else begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:543:7
			norm_shamt = addend_shamt_q;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:544:7
			normalized_exponent = tentative_exponent_q;
		end
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:549:3
	assign sum_shifted = sum_q << norm_shamt;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:553:3
	always @(*) begin : small_norm
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:555:5
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:556:5
		final_exponent = normalized_exponent;
		// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:559:5
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:560:7
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:561:7
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:567:7
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:568:7
			final_exponent = normalized_exponent - 1;
		end
		else
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:571:7
			final_exponent = 1'sb0;
	end
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:576:3
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:581:3
	wire pre_round_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:582:3
	wire [EXP_BITS - 1:0] pre_round_exponent;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:583:3
	wire [MAN_BITS - 1:0] pre_round_mantissa;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:584:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] pre_round_abs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:585:3
	wire [1:0] round_sticky_bits;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:587:3
	wire of_before_round;
	wire of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:588:3
	wire uf_before_round;
	wire uf_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:589:3
	wire result_zero;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:591:3
	wire rounded_sign;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:592:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] rounded_abs;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:595:3
	assign of_before_round = final_exponent >= ((2 ** EXP_BITS) - 1);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:596:3
	assign uf_before_round = final_exponent == 0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:599:3
	assign pre_round_sign = final_sign_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:600:3
	assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : $unsigned(final_exponent[EXP_BITS - 1:0]));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:601:3
	assign pre_round_mantissa = (of_before_round ? {MAN_BITS {1'sb1}} : final_mantissa[MAN_BITS:1]);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:602:3
	assign pre_round_abs = {pre_round_exponent, pre_round_mantissa};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:605:3
	assign round_sticky_bits = (of_before_round ? 2'b11 : {final_mantissa[0], sticky_after_norm});
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:608:3
	fpnew_rounding #(.AbsWidth(EXP_BITS + MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:622:3
	assign uf_after_round = (rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}}) || (((pre_round_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}}) && (rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == 1)) && ((round_sticky_bits != 2'b11) || (!sum_sticky_bits[(MAN_BITS * 2) + 4] && ((rnd_mode_q == 3'b000) || (rnd_mode_q == 3'b100)))));
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:625:3
	assign of_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:630:3
	wire [WIDTH - 1:0] regular_result;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:631:3
	wire [4:0] regular_status;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:634:3
	assign regular_result = {rounded_sign, rounded_abs};
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:635:3
	assign regular_status[4] = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:636:3
	assign regular_status[3] = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:637:3
	assign regular_status[2] = of_before_round | of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:638:3
	assign regular_status[1] = uf_after_round & regular_status[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:639:3
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:642:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:643:3
	wire [4:0] status_d;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:646:3
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:647:3
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:653:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:654:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:655:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) - 1)) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))) + (TagType_TagType_TagType_TagType_TAG_WIDTH - 1))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAG_WIDTH + 1) : (TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))) : ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] out_pipe_tag_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:656:3
	reg [0:NUM_OUT_REGS] out_pipe_mask_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:657:3
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:658:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:660:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:663:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_0252C;
	assign sv2v_tmp_0252C = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_0252C;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:664:3
	wire [5:1] sv2v_tmp_2A843;
	assign sv2v_tmp_2A843 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_2A843;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:665:3
	wire [((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)) * 1:1] sv2v_tmp_46F05;
	assign sv2v_tmp_46F05 = mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_tmp_46F05;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:666:3
	wire [1:1] sv2v_tmp_DB780;
	assign sv2v_tmp_DB780 = mid_pipe_mask_q[NUM_MID_REGS];
	always @(*) out_pipe_mask_q[0] = sv2v_tmp_DB780;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:667:3
	wire [1:1] sv2v_tmp_9E262;
	assign sv2v_tmp_9E262 = mid_pipe_aux_q[NUM_MID_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_9E262;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:668:3
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:670:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:672:3
	genvar _gv_i_235;
	generate
		for (_gv_i_235 = 0; _gv_i_235 < NUM_OUT_REGS; _gv_i_235 = _gv_i_235 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_235;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:674:5
			wire reg_ena;
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:678:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:680:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:680:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:680:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at /vortex/third_party/cvfpu/src/fpnew_fma.sv:680:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:682:5
			assign reg_ena = (out_pipe_ready[i] & out_pipe_valid_q[i]) | reg_ena_i[(NUM_INP_REGS + NUM_MID_REGS) + i];
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:684:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:684:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:684:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:684:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:685:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:685:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:685:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:685:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:686:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:686:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:686:189
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= sv2v_cast_48BE4(1'sb0);
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:686:297
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:687:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:687:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:687:179
					out_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:687:287
					out_pipe_mask_q[i + 1] <= (reg_ena ? out_pipe_mask_q[i] : out_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:688:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:688:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:688:189
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at /vortex/third_party/cvfpu/src/fpnew_fma.sv:688:297
					out_pipe_aux_q[i + 1] <= (reg_ena ? out_pipe_aux_q[i] : out_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:691:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:693:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:694:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:695:3
	assign extension_bit_o = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:696:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAG_WIDTH + 0) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0)))+:((TagType_TagType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? TagType_TagType_TagType_TagType_TAG_WIDTH + 1 : 1 - (TagType_TagType_TagType_TagType_TAG_WIDTH + 0))];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:697:3
	assign mask_o = out_pipe_mask_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:698:3
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:699:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: /vortex/third_party/cvfpu/src/fpnew_fma.sv:700:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
// removed package "cb_filter_pkg"
// removed interface: STREAM_DV
module rr_arb_tree_4016C_91833 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	req_o,
	gnt_i,
	data_o,
	idx_o
);
	// removed localparam type DataType_TagType_TagType_TAG_WIDTH_type
	// removed localparam type DataType_Width_type
	parameter signed [31:0] DataType_TagType_TagType_TAG_WIDTH = 0;
	parameter [31:0] DataType_Width = 0;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:49:13
	parameter [31:0] NumIn = 64;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:51:13
	parameter [31:0] DataWidth = 32;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:53:26
	// removed localparam type DataType
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:60:13
	parameter [0:0] ExtPrio = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:67:13
	parameter [0:0] AxiVldRdy = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:74:13
	parameter [0:0] LockIn = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:78:13
	parameter [0:0] FairArb = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:81:13
	parameter [31:0] IdxWidth = (NumIn > 32'd1 ? $unsigned($clog2(NumIn)) : 32'd1);
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:84:26
	// removed localparam type idx_t
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:87:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:89:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:91:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:93:3
	input wire [IdxWidth - 1:0] rr_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:95:3
	input wire [NumIn - 1:0] req_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:98:3
	output wire [NumIn - 1:0] gnt_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:101:3
	input wire [(NumIn * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))) - 1:0] data_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:103:3
	output wire req_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:105:3
	input wire gnt_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:107:3
	output wire [((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))) - 1:0] data_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:109:3
	output wire [IdxWidth - 1:0] idx_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:122:3
	function automatic [IdxWidth - 1:0] sv2v_cast_29535;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_29535 = inp;
	endfunction
	function automatic [((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))) - 1:0] sv2v_cast_790D3;
		input reg [((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))) - 1:0] inp;
		sv2v_cast_790D3 = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : gen_pass_through
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:123:5
			assign req_o = req_i[0];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:124:5
			assign gnt_o[0] = gnt_i;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:125:5
			assign data_o = data_i[0+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:126:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_arbiter
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:129:5
			localparam [31:0] NumLevels = $unsigned($clog2(NumIn));
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:132:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * IdxWidth) - 1 : ((3 - (2 ** NumLevels)) * IdxWidth) + ((((2 ** NumLevels) - 2) * IdxWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * IdxWidth)] index_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:133:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))) - 1 : ((3 - (2 ** NumLevels)) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))) + ((((2 ** NumLevels) - 2) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))))] data_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:134:5
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:135:5
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:137:5
			reg [IdxWidth - 1:0] rr_q;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:138:5
			wire [NumIn - 1:0] req_d;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:141:5
			assign req_o = req_nodes[0];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:142:5
			assign data_o = data_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:143:5
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * IdxWidth+:IdxWidth];
			if (ExtPrio) begin : gen_ext_rr
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:146:7
				wire [IdxWidth:1] sv2v_tmp_4C2F0;
				assign sv2v_tmp_4C2F0 = rr_i;
				always @(*) rr_q = sv2v_tmp_4C2F0;
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:147:7
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:149:7
				wire [IdxWidth - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:153:9
					wire lock_d;
					reg lock_q;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:154:9
					reg [NumIn - 1:0] req_q;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:156:9
					assign lock_d = req_o & ~gnt_i;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:157:9
					assign req_d = (lock_q ? req_q : req_i);
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:159:9
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:160:11
						if (!rst_ni)
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:161:13
							lock_q <= 1'sb0;
						else
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:163:13
							if (flush_i)
								// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:164:15
								lock_q <= 1'sb0;
							else
								// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:166:15
								lock_q <= lock_d;
					end
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:173:11
					// removed an assertion item
					// lock : assert property (@(posedge clk_i) 
					// 	(LockIn |-> (req_o && !gnt_i |=> idx_o == $past(idx_o)))
					// ) else begin
					// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:175:17
					// 	$fatal(1, "Lock implies same arbiter decision in next cycle if output is not                             ready.");
					// end
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:178:11
					wire [NumIn - 1:0] req_tmp;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:179:11
					assign req_tmp = req_q & req_i;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:180:11
					// removed an assertion item
					// lock_req : assume property (@(posedge clk_i) 
					// 	(LockIn |-> (lock_d |=> req_tmp == req_q))
					// ) else begin
					// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:182:17
					// 	$fatal(1, "It is disallowed to deassert unserved request signals when LockIn is                             enabled.");
					// end
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:187:9
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:188:11
						if (!rst_ni)
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:189:13
							req_q <= 1'sb0;
						else
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:191:13
							if (flush_i)
								// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:192:15
								req_q <= 1'sb0;
							else
								// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:194:15
								req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:199:9
					assign req_d = req_i;
				end
				if (FairArb) begin : gen_fair_arb
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:203:9
					wire [NumIn - 1:0] upper_mask;
					wire [NumIn - 1:0] lower_mask;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:204:9
					wire [IdxWidth - 1:0] upper_idx;
					wire [IdxWidth - 1:0] lower_idx;
					wire [IdxWidth - 1:0] next_idx;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:205:9
					wire upper_empty;
					wire lower_empty;
					genvar _gv_i_251;
					for (_gv_i_251 = 0; _gv_i_251 < NumIn; _gv_i_251 = _gv_i_251 + 1) begin : gen_mask
						localparam i = _gv_i_251;
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:208:11
						assign upper_mask[i] = (i > rr_q ? req_d[i] : 1'b0);
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:209:11
						assign lower_mask[i] = (i <= rr_q ? req_d[i] : 1'b0);
					end
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:212:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_upper(
						.in_i(upper_mask),
						.cnt_o(upper_idx),
						.empty_o(upper_empty)
					);
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:221:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_lower(
						.in_i(lower_mask),
						.cnt_o(lower_idx),
						.empty_o()
					);
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:230:9
					assign next_idx = (upper_empty ? lower_idx : upper_idx);
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:231:9
					assign rr_d = (gnt_i && req_o ? next_idx : rr_q);
				end
				else begin : gen_unfair_arb
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:234:9
					assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_29535(NumIn - 1) ? {IdxWidth {1'sb0}} : rr_q + 1'b1) : rr_q);
				end
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:238:7
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:239:9
					if (!rst_ni)
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:240:11
						rr_q <= 1'sb0;
					else
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:242:11
						if (flush_i)
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:243:13
							rr_q <= 1'sb0;
						else
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:245:13
							rr_q <= rr_d;
				end
			end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:251:5
			assign gnt_nodes[0] = gnt_i;
			genvar _gv_level_1;
			for (_gv_level_1 = 0; $unsigned(_gv_level_1) < NumLevels; _gv_level_1 = _gv_level_1 + 1) begin : gen_levels
				localparam level = _gv_level_1;
				genvar _gv_l_1;
				for (_gv_l_1 = 0; _gv_l_1 < (2 ** level); _gv_l_1 = _gv_l_1 + 1) begin : gen_level
					localparam l = _gv_l_1;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:257:9
					wire sel;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:259:9
					localparam [31:0] Idx0 = ((2 ** level) - 1) + l;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:260:9
					localparam [31:0] Idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : gen_reduce
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:266:13
							assign req_nodes[Idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:269:13
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:271:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_29535(sel);
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:272:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))] = (sel ? data_i[((l * 2) + 1) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))] : data_i[(l * 2) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))]);
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:273:13
							assign gnt_o[l * 2] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:274:13
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : gen_first
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:278:13
							assign req_nodes[Idx0] = req_d[l * 2];
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:279:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = 1'sb0;
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:280:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))] = data_i[(l * 2) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))];
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:281:13
							assign gnt_o[l * 2] = gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : gen_out_of_range
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:285:13
							assign req_nodes[Idx0] = 1'b0;
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:286:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_29535(1'sb0);
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:287:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))] = sv2v_cast_790D3(1'sb0);
						end
					end
					else begin : gen_other_levels
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:292:11
						assign req_nodes[Idx0] = req_nodes[Idx1] | req_nodes[Idx1 + 1];
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:295:11
						assign sel = ~req_nodes[Idx1] | (req_nodes[Idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:297:11
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = (sel ? sv2v_cast_29535({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_29535({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:301:11
						assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))] = (sel ? data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))] : data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * ((DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0)))+:(DataType_Width + 6) + ((DataType_TagType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TagType_TAG_WIDTH + 0))]);
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:302:11
						assign gnt_nodes[Idx1] = gnt_nodes[Idx0] & ~sel;
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:303:11
						assign gnt_nodes[Idx1 + 1] = gnt_nodes[Idx0] & sel;
					end
				end
			end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:312:5
			initial begin : p_assert
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:313:7
			end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:319:5
			// removed an assertion item
			// hot_one : assert property (@(posedge clk_i) 
			// 	$onehot0(gnt_o)
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:321:14
			// 	$fatal(1, "Grant signal must be hot1 or zero.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:323:5
			// removed an assertion item
			// gnt0 : assert property (@(posedge clk_i) 
			// 	(|gnt_o |-> gnt_i)
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:325:14
			// 	$fatal(1, "Grant out implies grant in.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:327:5
			// removed an assertion item
			// gnt1 : assert property (@(posedge clk_i) 
			// 	(req_o |-> (gnt_i |-> |gnt_o))
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:329:14
			// 	$fatal(1, "Req out and grant in implies grant out.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:331:5
			// removed an assertion item
			// gnt_idx : assert property (@(posedge clk_i) 
			// 	(req_o |-> (gnt_i |-> gnt_o[idx_o]))
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:333:14
			// 	$fatal(1, "Idx_o / gnt_o do not match.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:335:5
			// removed an assertion item
			// req0 : assert property (@(posedge clk_i) 
			// 	(|req_i |-> req_o)
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:337:14
			// 	$fatal(1, "Req in implies req out.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:339:5
			// removed an assertion item
			// req1 : assert property (@(posedge clk_i) 
			// 	(req_o |-> |req_i)
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:341:14
			// 	$fatal(1, "Req out implies req in.");
			// end
		end
	endgenerate
endmodule
module rr_arb_tree_CF21D_98F90 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	req_o,
	gnt_i,
	data_o,
	idx_o
);
	// removed localparam type DataType_TagType_TAG_WIDTH_type
	// removed localparam type DataType_WIDTH_type
	parameter signed [31:0] DataType_TagType_TAG_WIDTH = 0;
	parameter [31:0] DataType_WIDTH = 0;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:49:13
	parameter [31:0] NumIn = 64;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:51:13
	parameter [31:0] DataWidth = 32;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:53:26
	// removed localparam type DataType
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:60:13
	parameter [0:0] ExtPrio = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:67:13
	parameter [0:0] AxiVldRdy = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:74:13
	parameter [0:0] LockIn = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:78:13
	parameter [0:0] FairArb = 1'b1;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:81:13
	parameter [31:0] IdxWidth = (NumIn > 32'd1 ? $unsigned($clog2(NumIn)) : 32'd1);
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:84:26
	// removed localparam type idx_t
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:87:3
	input wire clk_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:89:3
	input wire rst_ni;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:91:3
	input wire flush_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:93:3
	input wire [IdxWidth - 1:0] rr_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:95:3
	input wire [NumIn - 1:0] req_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:98:3
	output wire [NumIn - 1:0] gnt_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:101:3
	input wire [(NumIn * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))) - 1:0] data_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:103:3
	output wire req_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:105:3
	input wire gnt_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:107:3
	output wire [((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))) - 1:0] data_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:109:3
	output wire [IdxWidth - 1:0] idx_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:122:3
	function automatic [IdxWidth - 1:0] sv2v_cast_29535;
		input reg [IdxWidth - 1:0] inp;
		sv2v_cast_29535 = inp;
	endfunction
	function automatic [((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))) - 1:0] sv2v_cast_7CC9D;
		input reg [((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))) - 1:0] inp;
		sv2v_cast_7CC9D = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : gen_pass_through
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:123:5
			assign req_o = req_i[0];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:124:5
			assign gnt_o[0] = gnt_i;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:125:5
			assign data_o = data_i[0+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:126:5
			assign idx_o = 1'sb0;
		end
		else begin : gen_arbiter
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:129:5
			localparam [31:0] NumLevels = $unsigned($clog2(NumIn));
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:132:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * IdxWidth) - 1 : ((3 - (2 ** NumLevels)) * IdxWidth) + ((((2 ** NumLevels) - 2) * IdxWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * IdxWidth)] index_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:133:5
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))) - 1 : ((3 - (2 ** NumLevels)) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))) + ((((2 ** NumLevels) - 2) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))))] data_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:134:5
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:135:5
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:137:5
			reg [IdxWidth - 1:0] rr_q;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:138:5
			wire [NumIn - 1:0] req_d;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:141:5
			assign req_o = req_nodes[0];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:142:5
			assign data_o = data_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:143:5
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * IdxWidth+:IdxWidth];
			if (ExtPrio) begin : gen_ext_rr
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:146:7
				wire [IdxWidth:1] sv2v_tmp_4C2F0;
				assign sv2v_tmp_4C2F0 = rr_i;
				always @(*) rr_q = sv2v_tmp_4C2F0;
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:147:7
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:149:7
				wire [IdxWidth - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:153:9
					wire lock_d;
					reg lock_q;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:154:9
					reg [NumIn - 1:0] req_q;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:156:9
					assign lock_d = req_o & ~gnt_i;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:157:9
					assign req_d = (lock_q ? req_q : req_i);
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:159:9
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:160:11
						if (!rst_ni)
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:161:13
							lock_q <= 1'sb0;
						else
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:163:13
							if (flush_i)
								// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:164:15
								lock_q <= 1'sb0;
							else
								// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:166:15
								lock_q <= lock_d;
					end
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:173:11
					// removed an assertion item
					// lock : assert property (@(posedge clk_i) 
					// 	(LockIn |-> (req_o && !gnt_i |=> idx_o == $past(idx_o)))
					// ) else begin
					// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:175:17
					// 	$fatal(1, "Lock implies same arbiter decision in next cycle if output is not                             ready.");
					// end
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:178:11
					wire [NumIn - 1:0] req_tmp;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:179:11
					assign req_tmp = req_q & req_i;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:180:11
					// removed an assertion item
					// lock_req : assume property (@(posedge clk_i) 
					// 	(LockIn |-> (lock_d |=> req_tmp == req_q))
					// ) else begin
					// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:182:17
					// 	$fatal(1, "It is disallowed to deassert unserved request signals when LockIn is                             enabled.");
					// end
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:187:9
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:188:11
						if (!rst_ni)
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:189:13
							req_q <= 1'sb0;
						else
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:191:13
							if (flush_i)
								// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:192:15
								req_q <= 1'sb0;
							else
								// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:194:15
								req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:199:9
					assign req_d = req_i;
				end
				if (FairArb) begin : gen_fair_arb
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:203:9
					wire [NumIn - 1:0] upper_mask;
					wire [NumIn - 1:0] lower_mask;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:204:9
					wire [IdxWidth - 1:0] upper_idx;
					wire [IdxWidth - 1:0] lower_idx;
					wire [IdxWidth - 1:0] next_idx;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:205:9
					wire upper_empty;
					wire lower_empty;
					genvar _gv_i_251;
					for (_gv_i_251 = 0; _gv_i_251 < NumIn; _gv_i_251 = _gv_i_251 + 1) begin : gen_mask
						localparam i = _gv_i_251;
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:208:11
						assign upper_mask[i] = (i > rr_q ? req_d[i] : 1'b0);
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:209:11
						assign lower_mask[i] = (i <= rr_q ? req_d[i] : 1'b0);
					end
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:212:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_upper(
						.in_i(upper_mask),
						.cnt_o(upper_idx),
						.empty_o(upper_empty)
					);
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:221:9
					lzc #(
						.WIDTH(NumIn),
						.MODE(1'b0)
					) i_lzc_lower(
						.in_i(lower_mask),
						.cnt_o(lower_idx),
						.empty_o()
					);
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:230:9
					assign next_idx = (upper_empty ? lower_idx : upper_idx);
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:231:9
					assign rr_d = (gnt_i && req_o ? next_idx : rr_q);
				end
				else begin : gen_unfair_arb
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:234:9
					assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_29535(NumIn - 1) ? {IdxWidth {1'sb0}} : rr_q + 1'b1) : rr_q);
				end
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:238:7
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:239:9
					if (!rst_ni)
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:240:11
						rr_q <= 1'sb0;
					else
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:242:11
						if (flush_i)
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:243:13
							rr_q <= 1'sb0;
						else
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:245:13
							rr_q <= rr_d;
				end
			end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:251:5
			assign gnt_nodes[0] = gnt_i;
			genvar _gv_level_1;
			for (_gv_level_1 = 0; $unsigned(_gv_level_1) < NumLevels; _gv_level_1 = _gv_level_1 + 1) begin : gen_levels
				localparam level = _gv_level_1;
				genvar _gv_l_1;
				for (_gv_l_1 = 0; _gv_l_1 < (2 ** level); _gv_l_1 = _gv_l_1 + 1) begin : gen_level
					localparam l = _gv_l_1;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:257:9
					wire sel;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:259:9
					localparam [31:0] Idx0 = ((2 ** level) - 1) + l;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:260:9
					localparam [31:0] Idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : gen_reduce
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:266:13
							assign req_nodes[Idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:269:13
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:271:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_29535(sel);
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:272:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))] = (sel ? data_i[((l * 2) + 1) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))] : data_i[(l * 2) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))]);
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:273:13
							assign gnt_o[l * 2] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:274:13
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[Idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : gen_first
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:278:13
							assign req_nodes[Idx0] = req_d[l * 2];
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:279:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = 1'sb0;
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:280:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))] = data_i[(l * 2) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))];
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:281:13
							assign gnt_o[l * 2] = gnt_nodes[Idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : gen_out_of_range
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:285:13
							assign req_nodes[Idx0] = 1'b0;
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:286:13
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = sv2v_cast_29535(1'sb0);
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:287:13
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))] = sv2v_cast_7CC9D(1'sb0);
						end
					end
					else begin : gen_other_levels
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:292:11
						assign req_nodes[Idx0] = req_nodes[Idx1] | req_nodes[Idx1 + 1];
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:295:11
						assign sel = ~req_nodes[Idx1] | (req_nodes[Idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:297:11
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * IdxWidth+:IdxWidth] = (sel ? sv2v_cast_29535({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_29535({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * IdxWidth) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:301:11
						assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx0 : ((2 ** NumLevels) - 2) - Idx0) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))] = (sel ? data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 + 1 : ((2 ** NumLevels) - 2) - (Idx1 + 1)) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))] : data_nodes[(((2 ** NumLevels) - 2) >= 0 ? Idx1 : ((2 ** NumLevels) - 2) - Idx1) * ((DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0)))+:(DataType_WIDTH + 5) + ((DataType_TagType_TAG_WIDTH + 0) >= 0 ? DataType_TagType_TAG_WIDTH + 1 : 1 - (DataType_TagType_TAG_WIDTH + 0))]);
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:302:11
						assign gnt_nodes[Idx1] = gnt_nodes[Idx0] & ~sel;
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:303:11
						assign gnt_nodes[Idx1 + 1] = gnt_nodes[Idx0] & sel;
					end
				end
			end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:312:5
			initial begin : p_assert
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:313:7
			end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:319:5
			// removed an assertion item
			// hot_one : assert property (@(posedge clk_i) 
			// 	$onehot0(gnt_o)
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:321:14
			// 	$fatal(1, "Grant signal must be hot1 or zero.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:323:5
			// removed an assertion item
			// gnt0 : assert property (@(posedge clk_i) 
			// 	(|gnt_o |-> gnt_i)
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:325:14
			// 	$fatal(1, "Grant out implies grant in.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:327:5
			// removed an assertion item
			// gnt1 : assert property (@(posedge clk_i) 
			// 	(req_o |-> (gnt_i |-> |gnt_o))
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:329:14
			// 	$fatal(1, "Req out and grant in implies grant out.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:331:5
			// removed an assertion item
			// gnt_idx : assert property (@(posedge clk_i) 
			// 	(req_o |-> (gnt_i |-> gnt_o[idx_o]))
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:333:14
			// 	$fatal(1, "Idx_o / gnt_o do not match.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:335:5
			// removed an assertion item
			// req0 : assert property (@(posedge clk_i) 
			// 	(|req_i |-> req_o)
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:337:14
			// 	$fatal(1, "Req in implies req out.");
			// end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:339:5
			// removed an assertion item
			// req1 : assert property (@(posedge clk_i) 
			// 	(req_o |-> |req_i)
			// ) else begin
			// 	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/rr_arb_tree.sv:341:14
			// 	$fatal(1, "Req out implies req in.");
			// end
		end
	endgenerate
endmodule
// removed package "cf_math_pkg"
module popcount (
	data_i,
	popcount_o
);
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:20:15
	parameter [31:0] INPUT_WIDTH = 256;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:21:16
	localparam [31:0] PopcountWidth = $clog2(INPUT_WIDTH) + 1;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:23:5
	input wire [INPUT_WIDTH - 1:0] data_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:24:5
	output wire [PopcountWidth - 1:0] popcount_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:27:4
	localparam [31:0] PaddedWidth = 1 << $clog2(INPUT_WIDTH);
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:29:4
	reg [PaddedWidth - 1:0] padded_input;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:30:4
	wire [PopcountWidth - 2:0] left_child_result;
	wire [PopcountWidth - 2:0] right_child_result;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:33:4
	always @(*) begin
		// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:34:6
		padded_input = 1'sb0;
		// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:35:6
		padded_input[INPUT_WIDTH - 1:0] = data_i;
	end
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:39:4
	generate
		if (INPUT_WIDTH == 1) begin : single_node
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:40:6
			assign left_child_result = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:41:6
			assign right_child_result = padded_input[0];
		end
		else if (INPUT_WIDTH == 2) begin : leaf_node
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:43:6
			assign left_child_result = padded_input[1];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:44:6
			assign right_child_result = padded_input[0];
		end
		else begin : non_leaf_node
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:46:6
			popcount #(.INPUT_WIDTH(PaddedWidth / 2)) left_child(
				.data_i(padded_input[PaddedWidth - 1:PaddedWidth / 2]),
				.popcount_o(left_child_result)
			);
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:51:6
			popcount #(.INPUT_WIDTH(PaddedWidth / 2)) right_child(
				.data_i(padded_input[(PaddedWidth / 2) - 1:0]),
				.popcount_o(right_child_result)
			);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/popcount.sv:58:4
	assign popcount_o = left_child_result + right_child_result;
endmodule
// removed package "ecc_pkg"
module lzc (
	in_i,
	cnt_o,
	empty_o
);
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:27:13
	parameter [31:0] WIDTH = 2;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:29:13
	parameter [0:0] MODE = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:33:13
	function automatic [31:0] cf_math_pkg_idx_width;
		// Trace: /vortex/third_party/cvfpu/src/common_cells/src/cf_math_pkg.sv:57:52
		input reg [31:0] num_idx;
		// Trace: /vortex/third_party/cvfpu/src/common_cells/src/cf_math_pkg.sv:58:9
		cf_math_pkg_idx_width = (num_idx > 32'd1 ? $unsigned($clog2(num_idx)) : 32'd1);
	endfunction
	parameter [31:0] CNT_WIDTH = cf_math_pkg_idx_width(WIDTH);
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:36:3
	input wire [WIDTH - 1:0] in_i;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:38:3
	output wire [CNT_WIDTH - 1:0] cnt_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:40:3
	output wire empty_o;
	// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:43:3
	generate
		if (WIDTH == 1) begin : gen_degenerate_lzc
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:45:5
			assign cnt_o[0] = !in_i[0];
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:46:5
			assign empty_o = !in_i[0];
		end
		else begin : gen_lzc
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:50:5
			localparam [31:0] NumLevels = $clog2(WIDTH);
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:53:5
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:58:5
			wire [(WIDTH * NumLevels) - 1:0] index_lut;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:59:5
			wire [(2 ** NumLevels) - 1:0] sel_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:60:5
			wire [((2 ** NumLevels) * NumLevels) - 1:0] index_nodes;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:62:5
			reg [WIDTH - 1:0] in_tmp;
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:65:5
			always @(*) begin : flip_vector
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:66:7
				begin : sv2v_autoblock_1
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:66:12
					reg [31:0] i;
					// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:66:12
					for (i = 0; i < WIDTH; i = i + 1)
						begin
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:67:9
							in_tmp[i] = (MODE ? in_i[(WIDTH - 1) - i] : in_i[i]);
						end
				end
			end
			genvar _gv_j_29;
			for (_gv_j_29 = 0; $unsigned(_gv_j_29) < WIDTH; _gv_j_29 = _gv_j_29 + 1) begin : g_index_lut
				localparam j = _gv_j_29;
				// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:72:7
				function automatic [NumLevels - 1:0] sv2v_cast_5699A;
					input reg [NumLevels - 1:0] inp;
					sv2v_cast_5699A = inp;
				endfunction
				assign index_lut[j * NumLevels+:NumLevels] = sv2v_cast_5699A($unsigned(j));
			end
			genvar _gv_level_2;
			for (_gv_level_2 = 0; $unsigned(_gv_level_2) < NumLevels; _gv_level_2 = _gv_level_2 + 1) begin : g_levels
				localparam level = _gv_level_2;
				if ($unsigned(level) == (NumLevels - 1)) begin : g_last_level
					genvar _gv_k_4;
					for (_gv_k_4 = 0; _gv_k_4 < (2 ** level); _gv_k_4 = _gv_k_4 + 1) begin : g_level
						localparam k = _gv_k_4;
						if (($unsigned(k) * 2) < (WIDTH - 1)) begin : g_reduce
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:80:13
							assign sel_nodes[((2 ** level) - 1) + k] = in_tmp[k * 2] | in_tmp[(k * 2) + 1];
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:81:13
							assign index_nodes[(((2 ** level) - 1) + k) * NumLevels+:NumLevels] = (in_tmp[k * 2] == 1'b1 ? index_lut[(k * 2) * NumLevels+:NumLevels] : index_lut[((k * 2) + 1) * NumLevels+:NumLevels]);
						end
						if (($unsigned(k) * 2) == (WIDTH - 1)) begin : g_base
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:87:13
							assign sel_nodes[((2 ** level) - 1) + k] = in_tmp[k * 2];
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:88:13
							assign index_nodes[(((2 ** level) - 1) + k) * NumLevels+:NumLevels] = index_lut[(k * 2) * NumLevels+:NumLevels];
						end
						if (($unsigned(k) * 2) > (WIDTH - 1)) begin : g_out_of_range
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:92:13
							assign sel_nodes[((2 ** level) - 1) + k] = 1'b0;
							// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:93:13
							assign index_nodes[(((2 ** level) - 1) + k) * NumLevels+:NumLevels] = 1'sb0;
						end
					end
				end
				else begin : g_not_last_level
					genvar _gv_l_2;
					for (_gv_l_2 = 0; _gv_l_2 < (2 ** level); _gv_l_2 = _gv_l_2 + 1) begin : g_level
						localparam l = _gv_l_2;
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:98:11
						assign sel_nodes[((2 ** level) - 1) + l] = sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] | sel_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) + 1];
						// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:100:11
						assign index_nodes[(((2 ** level) - 1) + l) * NumLevels+:NumLevels] = (sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] == 1'b1 ? index_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) * NumLevels+:NumLevels] : index_nodes[((((2 ** (level + 1)) - 1) + (l * 2)) + 1) * NumLevels+:NumLevels]);
					end
				end
			end
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:107:5
			assign cnt_o = (NumLevels > $unsigned(0) ? index_nodes[0+:NumLevels] : {$clog2(WIDTH) {1'b0}});
			// Trace: /vortex/third_party/cvfpu/src/common_cells/src/lzc.sv:108:5
			assign empty_o = (NumLevels > $unsigned(0) ? ~sel_nodes[0] : ~(|in_i));
		end
	endgenerate
endmodule
// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:41:1
// removed ["import defs_div_sqrt_mvp::*;"]
module control_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Start_SI,
	Kill_SI,
	Special_case_SBI,
	Special_case_dly_SBI,
	Precision_ctl_SI,
	Format_sel_SI,
	Numerator_DI,
	Exp_num_DI,
	Denominator_DI,
	Exp_den_DI,
	Div_start_dly_SO,
	Sqrt_start_dly_SO,
	Div_enable_SO,
	Sqrt_enable_SO,
	Full_precision_SO,
	FP32_SO,
	FP64_SO,
	FP16_SO,
	FP16ALT_SO,
	Ready_SO,
	Done_SO,
	Mant_result_prenorm_DO,
	Exp_result_prenorm_DO
);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:46:4
	input wire Clk_CI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:47:4
	input wire Rst_RBI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:48:4
	input wire Div_start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:49:4
	input wire Sqrt_start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:50:4
	input wire Start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:51:4
	input wire Kill_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:52:4
	input wire Special_case_SBI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:53:4
	input wire Special_case_dly_SBI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:54:4
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:55:4
	input wire [1:0] Format_sel_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:56:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Numerator_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:57:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_num_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:58:4
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Denominator_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:59:4
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_den_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:62:4
	output wire Div_start_dly_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:63:4
	output wire Sqrt_start_dly_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:64:4
	output reg Div_enable_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:65:4
	output reg Sqrt_enable_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:69:4
	output wire Full_precision_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:70:4
	output wire FP32_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:71:4
	output wire FP64_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:72:4
	output wire FP16_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:73:4
	output wire FP16ALT_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:75:4
	output reg Ready_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:76:4
	output reg Done_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:78:4
	output reg [56:0] Mant_result_prenorm_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:80:4
	output wire [12:0] Exp_result_prenorm_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:83:4
	reg [57:0] Partial_remainder_DN;
	reg [57:0] Partial_remainder_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:84:4
	reg [56:0] Quotient_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:88:4
	wire [53:0] Numerator_se_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:89:4
	wire [53:0] Denominator_se_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:90:4
	reg [53:0] Denominator_se_DB;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:92:4
	assign Numerator_se_D = {1'b0, Numerator_DI};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:94:4
	assign Denominator_se_D = {1'b0, Denominator_DI};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:96:3
	localparam defs_div_sqrt_mvp_C_MANT_FP16 = 10;
	localparam defs_div_sqrt_mvp_C_MANT_FP16ALT = 7;
	localparam defs_div_sqrt_mvp_C_MANT_FP32 = 23;
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:98:6
		if (FP32_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:100:10
			Denominator_se_DB = {~Denominator_se_D[53:29], {29 {1'b0}}};
		else if (FP64_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:103:10
			Denominator_se_DB = ~Denominator_se_D;
		else if (FP16_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:106:10
			Denominator_se_DB = {~Denominator_se_D[53:42], {42 {1'b0}}};
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:109:10
			Denominator_se_DB = {~Denominator_se_D[53:45], {45 {1'b0}}};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:114:4
	wire [53:0] Mant_D_sqrt_Norm;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:116:4
	assign Mant_D_sqrt_Norm = (Exp_num_DI[0] ? {1'b0, Numerator_DI} : {Numerator_DI, 1'b0});
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:121:4
	reg [1:0] Format_sel_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:123:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:125:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:127:13
			Format_sel_S <= 'b0;
		else if (Start_SI && Ready_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:131:13
			Format_sel_S <= Format_sel_SI;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:135:13
			Format_sel_S <= Format_sel_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:139:4
	assign FP32_SO = Format_sel_S == 2'b00;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:140:4
	assign FP64_SO = Format_sel_S == 2'b01;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:141:4
	assign FP16_SO = Format_sel_S == 2'b10;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:142:4
	assign FP16ALT_SO = Format_sel_S == 2'b11;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:150:4
	reg [5:0] Precision_ctl_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:151:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:153:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:155:13
			Precision_ctl_S <= 'b0;
		else if (Start_SI && Ready_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:159:13
			Precision_ctl_S <= Precision_ctl_SI;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:163:13
			Precision_ctl_S <= Precision_ctl_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:166:3
	assign Full_precision_SO = Precision_ctl_S == 6'h00;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:170:6
	reg [5:0] State_ctl_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:171:6
	wire [5:0] State_Two_iteration_unit_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:172:6
	wire [5:0] State_Four_iteration_unit_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:174:5
	assign State_Two_iteration_unit_S = Precision_ctl_S[5:1];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:175:5
	assign State_Four_iteration_unit_S = Precision_ctl_S[5:2];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:176:6
	localparam defs_div_sqrt_mvp_Iteration_unit_num_S = 2'b10;
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:178:10
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:182:16
				case (Format_sel_S)
					2'b00:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:185:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:187:26
							State_ctl_S = 6'h1b;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:191:26
							State_ctl_S = Precision_ctl_S;
					2'b01:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:196:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:198:26
							State_ctl_S = 6'h38;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:202:26
							State_ctl_S = Precision_ctl_S;
					2'b10:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:207:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:209:26
							State_ctl_S = 6'h0e;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:213:26
							State_ctl_S = Precision_ctl_S;
					2'b11:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:218:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:220:26
							State_ctl_S = 6'h0b;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:224:26
							State_ctl_S = Precision_ctl_S;
				endcase
			2'b01:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:234:16
				case (Format_sel_S)
					2'b00:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:237:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:239:26
							State_ctl_S = 6'h0d;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:243:26
							State_ctl_S = State_Two_iteration_unit_S;
					2'b01:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:248:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:250:26
							State_ctl_S = 6'h1b;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:254:26
							State_ctl_S = State_Two_iteration_unit_S;
					2'b10:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:259:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:261:26
							State_ctl_S = 6'h06;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:265:26
							State_ctl_S = State_Two_iteration_unit_S;
					2'b11:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:270:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:272:26
							State_ctl_S = 6'h05;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:276:26
							State_ctl_S = State_Two_iteration_unit_S;
				endcase
			2'b10:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:286:16
				case (Format_sel_S)
					2'b00:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:289:22
						case (Precision_ctl_S)
							6'h00:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:292:28
								State_ctl_S = 6'h08;
							6'h06, 6'h07, 6'h08:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:296:28
								State_ctl_S = 6'h02;
							6'h09, 6'h0a, 6'h0b:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:300:28
								State_ctl_S = 6'h03;
							6'h0c, 6'h0d, 6'h0e:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:304:28
								State_ctl_S = 6'h04;
							6'h0f, 6'h10, 6'h11:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:308:28
								State_ctl_S = 6'h05;
							6'h12, 6'h13, 6'h14:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:312:28
								State_ctl_S = 6'h06;
							6'h15, 6'h16, 6'h17:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:316:28
								State_ctl_S = 6'h07;
							default:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:320:28
								State_ctl_S = 6'h08;
						endcase
					2'b01:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:326:22
						case (Precision_ctl_S)
							6'h00:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:329:28
								State_ctl_S = 6'h12;
							6'h06, 6'h07, 6'h08:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:333:28
								State_ctl_S = 6'h02;
							6'h09, 6'h0a, 6'h0b:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:337:28
								State_ctl_S = 6'h03;
							6'h0c, 6'h0d, 6'h0e:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:341:28
								State_ctl_S = 6'h04;
							6'h0f, 6'h10, 6'h11:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:345:28
								State_ctl_S = 6'h05;
							6'h12, 6'h13, 6'h14:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:349:28
								State_ctl_S = 6'h06;
							6'h15, 6'h16, 6'h17:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:353:28
								State_ctl_S = 6'h07;
							6'h18, 6'h19, 6'h1a:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:357:28
								State_ctl_S = 6'h08;
							6'h1b, 6'h1c, 6'h1d:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:361:28
								State_ctl_S = 6'h09;
							6'h1e, 6'h1f, 6'h20:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:365:28
								State_ctl_S = 6'h0a;
							6'h21, 6'h22, 6'h23:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:369:28
								State_ctl_S = 6'h0b;
							6'h24, 6'h25, 6'h26:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:373:28
								State_ctl_S = 6'h0c;
							6'h27, 6'h28, 6'h29:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:377:28
								State_ctl_S = 6'h0d;
							6'h2a, 6'h2b, 6'h2c:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:381:28
								State_ctl_S = 6'h0e;
							6'h2d, 6'h2e, 6'h2f:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:385:28
								State_ctl_S = 6'h0f;
							6'h30, 6'h31, 6'h32:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:389:28
								State_ctl_S = 6'h10;
							6'h33, 6'h34, 6'h35:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:393:28
								State_ctl_S = 6'h11;
							default:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:397:28
								State_ctl_S = 6'h12;
						endcase
					2'b10:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:403:22
						case (Precision_ctl_S)
							6'h00:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:406:28
								State_ctl_S = 6'h04;
							6'h06, 6'h07, 6'h08:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:410:28
								State_ctl_S = 6'h02;
							6'h09, 6'h0a, 6'h0b:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:414:28
								State_ctl_S = 6'h03;
							default:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:418:28
								State_ctl_S = 6'h04;
						endcase
					2'b11:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:424:22
						case (Precision_ctl_S)
							6'h00:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:427:28
								State_ctl_S = 6'h03;
							6'h06, 6'h07, 6'h08:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:431:28
								State_ctl_S = 6'h02;
							default:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:435:28
								State_ctl_S = 6'h03;
						endcase
				endcase
			2'b11:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:446:16
				case (Format_sel_S)
					2'b00:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:449:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:451:26
							State_ctl_S = 6'h06;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:455:26
							State_ctl_S = State_Four_iteration_unit_S;
					2'b01:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:460:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:462:26
							State_ctl_S = 6'h0d;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:466:26
							State_ctl_S = State_Four_iteration_unit_S;
					2'b10:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:471:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:473:26
							State_ctl_S = 6'h03;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:477:26
							State_ctl_S = State_Four_iteration_unit_S;
					2'b11:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:482:22
						if (Full_precision_SO)
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:484:26
							State_ctl_S = 6'h02;
						else
							// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:488:26
							State_ctl_S = State_Four_iteration_unit_S;
				endcase
		endcase
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:503:4
	reg Div_start_dly_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:505:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:507:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:509:13
			Div_start_dly_S <= 1'b0;
		else if (Div_start_SI && Ready_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:513:12
			Div_start_dly_S <= 1'b1;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:517:13
			Div_start_dly_S <= 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:521:4
	assign Div_start_dly_SO = Div_start_dly_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:523:3
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:524:5
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:525:7
			Div_enable_SO <= 1'b0;
		else if (Kill_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:528:7
			Div_enable_SO <= 1'b0;
		else if (Div_start_SI && Ready_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:530:7
			Div_enable_SO <= 1'b1;
		else if (Done_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:532:7
			Div_enable_SO <= 1'b0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:534:7
			Div_enable_SO <= Div_enable_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:537:4
	reg Sqrt_start_dly_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:539:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:541:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:543:13
			Sqrt_start_dly_S <= 1'b0;
		else if (Sqrt_start_SI && Ready_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:547:12
			Sqrt_start_dly_S <= 1'b1;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:551:13
			Sqrt_start_dly_S <= 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:554:5
	assign Sqrt_start_dly_SO = Sqrt_start_dly_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:556:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:557:5
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:558:7
			Sqrt_enable_SO <= 1'b0;
		else if (Kill_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:560:7
			Sqrt_enable_SO <= 1'b0;
		else if (Sqrt_start_SI && Ready_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:562:7
			Sqrt_enable_SO <= 1'b1;
		else if (Done_SO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:564:7
			Sqrt_enable_SO <= 1'b0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:566:7
			Sqrt_enable_SO <= Sqrt_enable_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:569:4
	reg [5:0] Crtl_cnt_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:570:4
	wire Start_dly_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:572:4
	assign Start_dly_S = Div_start_dly_S | Sqrt_start_dly_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:574:4
	wire Fsm_enable_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:575:4
	assign Fsm_enable_S = ((Start_dly_S | |Crtl_cnt_S) && ~Kill_SI) && Special_case_dly_SBI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:577:4
	wire Final_state_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:578:4
	assign Final_state_S = Crtl_cnt_S == State_ctl_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:581:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:583:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:585:14
			Crtl_cnt_S <= 1'sb0;
		else if (Final_state_S | Kill_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:589:15
			Crtl_cnt_S <= 1'sb0;
		else if (Fsm_enable_S)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:593:15
			Crtl_cnt_S <= Crtl_cnt_S + 1;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:597:15
			Crtl_cnt_S <= 1'sb0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:603:5
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:605:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:607:13
			Done_SO <= 1'b0;
		else if (Start_SI && Ready_SO) begin
			begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:611:13
				if (~Special_case_SBI)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:613:17
					Done_SO <= 1'b1;
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:617:17
					Done_SO <= 1'b0;
			end
		end
		else if (Final_state_S)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:622:13
			Done_SO <= 1'b1;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:626:13
			Done_SO <= 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:633:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:635:8
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:637:12
			Ready_SO <= 1'b1;
		else if (Start_SI && Ready_SO) begin
			begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:642:13
				if (~Special_case_SBI)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:644:17
					Ready_SO <= 1'b1;
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:648:17
					Ready_SO <= 1'b0;
			end
		end
		else if (Final_state_S | Kill_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:653:12
			Ready_SO <= 1'b1;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:657:12
			Ready_SO <= Ready_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:666:3
	wire Qcnt_one_0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:667:3
	wire Qcnt_one_1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:668:3
	wire [1:0] Qcnt_one_2;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:669:3
	wire [2:0] Qcnt_one_3;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:670:3
	wire [3:0] Qcnt_one_4;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:671:3
	wire [4:0] Qcnt_one_5;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:672:3
	wire [5:0] Qcnt_one_6;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:673:3
	wire [6:0] Qcnt_one_7;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:674:3
	wire [7:0] Qcnt_one_8;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:675:3
	wire [8:0] Qcnt_one_9;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:676:3
	wire [9:0] Qcnt_one_10;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:677:3
	wire [10:0] Qcnt_one_11;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:678:3
	wire [11:0] Qcnt_one_12;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:679:3
	wire [12:0] Qcnt_one_13;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:680:3
	wire [13:0] Qcnt_one_14;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:681:3
	wire [14:0] Qcnt_one_15;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:682:3
	wire [15:0] Qcnt_one_16;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:683:3
	wire [16:0] Qcnt_one_17;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:684:3
	wire [17:0] Qcnt_one_18;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:685:3
	wire [18:0] Qcnt_one_19;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:686:3
	wire [19:0] Qcnt_one_20;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:687:3
	wire [20:0] Qcnt_one_21;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:688:3
	wire [21:0] Qcnt_one_22;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:689:3
	wire [22:0] Qcnt_one_23;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:690:3
	wire [23:0] Qcnt_one_24;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:691:3
	wire [24:0] Qcnt_one_25;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:692:3
	wire [25:0] Qcnt_one_26;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:693:3
	wire [26:0] Qcnt_one_27;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:694:3
	wire [27:0] Qcnt_one_28;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:695:3
	wire [28:0] Qcnt_one_29;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:696:3
	wire [29:0] Qcnt_one_30;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:697:3
	wire [30:0] Qcnt_one_31;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:698:3
	wire [31:0] Qcnt_one_32;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:699:3
	wire [32:0] Qcnt_one_33;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:700:3
	wire [33:0] Qcnt_one_34;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:701:3
	wire [34:0] Qcnt_one_35;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:702:3
	wire [35:0] Qcnt_one_36;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:703:3
	wire [36:0] Qcnt_one_37;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:704:3
	wire [37:0] Qcnt_one_38;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:705:3
	wire [38:0] Qcnt_one_39;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:706:3
	wire [39:0] Qcnt_one_40;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:707:3
	wire [40:0] Qcnt_one_41;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:708:3
	wire [41:0] Qcnt_one_42;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:709:3
	wire [42:0] Qcnt_one_43;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:710:3
	wire [43:0] Qcnt_one_44;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:711:3
	wire [44:0] Qcnt_one_45;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:712:3
	wire [45:0] Qcnt_one_46;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:713:3
	wire [46:0] Qcnt_one_47;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:714:3
	wire [47:0] Qcnt_one_48;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:715:3
	wire [48:0] Qcnt_one_49;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:716:3
	wire [49:0] Qcnt_one_50;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:717:3
	wire [50:0] Qcnt_one_51;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:718:3
	wire [51:0] Qcnt_one_52;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:719:3
	wire [52:0] Qcnt_one_53;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:720:3
	wire [53:0] Qcnt_one_54;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:721:3
	wire [54:0] Qcnt_one_55;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:722:3
	wire [55:0] Qcnt_one_56;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:723:3
	wire [56:0] Qcnt_one_57;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:724:3
	wire [57:0] Qcnt_one_58;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:725:3
	wire [58:0] Qcnt_one_59;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:726:3
	wire [59:0] Qcnt_one_60;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:737:3
	wire [1:0] Qcnt_two_0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:738:3
	wire [2:0] Qcnt_two_1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:739:3
	wire [4:0] Qcnt_two_2;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:740:3
	wire [6:0] Qcnt_two_3;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:741:3
	wire [8:0] Qcnt_two_4;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:742:3
	wire [10:0] Qcnt_two_5;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:743:3
	wire [12:0] Qcnt_two_6;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:744:3
	wire [14:0] Qcnt_two_7;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:745:3
	wire [16:0] Qcnt_two_8;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:746:3
	wire [18:0] Qcnt_two_9;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:747:3
	wire [20:0] Qcnt_two_10;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:748:3
	wire [22:0] Qcnt_two_11;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:749:3
	wire [24:0] Qcnt_two_12;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:750:3
	wire [26:0] Qcnt_two_13;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:751:3
	wire [28:0] Qcnt_two_14;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:752:3
	wire [30:0] Qcnt_two_15;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:753:3
	wire [32:0] Qcnt_two_16;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:754:3
	wire [34:0] Qcnt_two_17;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:755:3
	wire [36:0] Qcnt_two_18;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:756:3
	wire [38:0] Qcnt_two_19;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:757:3
	wire [40:0] Qcnt_two_20;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:758:3
	wire [42:0] Qcnt_two_21;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:759:3
	wire [44:0] Qcnt_two_22;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:760:3
	wire [46:0] Qcnt_two_23;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:761:3
	wire [48:0] Qcnt_two_24;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:762:3
	wire [50:0] Qcnt_two_25;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:763:3
	wire [52:0] Qcnt_two_26;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:764:3
	wire [54:0] Qcnt_two_27;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:765:3
	wire [56:0] Qcnt_two_28;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:774:3
	wire [2:0] Qcnt_three_0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:775:3
	wire [4:0] Qcnt_three_1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:776:3
	wire [7:0] Qcnt_three_2;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:777:3
	wire [10:0] Qcnt_three_3;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:778:3
	wire [13:0] Qcnt_three_4;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:779:3
	wire [16:0] Qcnt_three_5;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:780:3
	wire [19:0] Qcnt_three_6;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:781:3
	wire [22:0] Qcnt_three_7;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:782:3
	wire [25:0] Qcnt_three_8;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:783:3
	wire [28:0] Qcnt_three_9;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:784:3
	wire [31:0] Qcnt_three_10;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:785:3
	wire [34:0] Qcnt_three_11;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:786:3
	wire [37:0] Qcnt_three_12;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:787:3
	wire [40:0] Qcnt_three_13;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:788:3
	wire [43:0] Qcnt_three_14;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:789:3
	wire [46:0] Qcnt_three_15;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:790:3
	wire [49:0] Qcnt_three_16;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:791:3
	wire [52:0] Qcnt_three_17;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:792:3
	wire [55:0] Qcnt_three_18;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:793:3
	wire [58:0] Qcnt_three_19;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:794:3
	wire [61:0] Qcnt_three_20;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:803:3
	wire [3:0] Qcnt_four_0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:804:3
	wire [6:0] Qcnt_four_1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:805:3
	wire [10:0] Qcnt_four_2;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:806:3
	wire [14:0] Qcnt_four_3;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:807:3
	wire [18:0] Qcnt_four_4;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:808:3
	wire [22:0] Qcnt_four_5;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:809:3
	wire [26:0] Qcnt_four_6;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:810:3
	wire [30:0] Qcnt_four_7;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:811:3
	wire [34:0] Qcnt_four_8;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:812:3
	wire [38:0] Qcnt_four_9;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:813:3
	wire [42:0] Qcnt_four_10;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:814:3
	wire [46:0] Qcnt_four_11;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:815:3
	wire [50:0] Qcnt_four_12;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:816:3
	wire [54:0] Qcnt_four_13;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:817:3
	wire [58:0] Qcnt_four_14;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:825:4
	wire [57:0] Sqrt_R0;
	reg [57:0] Sqrt_Q0;
	reg [57:0] Q_sqrt0;
	reg [57:0] Q_sqrt_com_0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:826:4
	wire [57:0] Sqrt_R1;
	reg [57:0] Sqrt_Q1;
	reg [57:0] Q_sqrt1;
	reg [57:0] Q_sqrt_com_1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:827:4
	wire [57:0] Sqrt_R2;
	reg [57:0] Sqrt_Q2;
	reg [57:0] Q_sqrt2;
	reg [57:0] Q_sqrt_com_2;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:828:4
	wire [57:0] Sqrt_R3;
	reg [57:0] Sqrt_Q3;
	reg [57:0] Q_sqrt3;
	reg [57:0] Q_sqrt_com_3;
	wire [57:0] Sqrt_R4;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:831:4
	reg [1:0] Sqrt_DI [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:832:4
	wire [1:0] Sqrt_DO [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:833:4
	wire Sqrt_carry_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:836:3
	wire [57:0] Iteration_cell_a_D [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:837:3
	wire [57:0] Iteration_cell_b_D [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:838:3
	wire [57:0] Iteration_cell_a_BMASK_D [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:839:3
	wire [57:0] Iteration_cell_b_BMASK_D [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:840:3
	wire Iteration_cell_carry_D [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:841:3
	wire [57:0] Iteration_cell_sum_D [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:842:3
	wire [57:0] Iteration_cell_sum_AMASK_D [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:845:3
	reg [3:0] Sqrt_quotinent_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:848:4
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:850:7
		case (Format_sel_S)
			2'b00: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:853:13
				Sqrt_quotinent_S = {~Iteration_cell_sum_AMASK_D[0][28], ~Iteration_cell_sum_AMASK_D[1][28], ~Iteration_cell_sum_AMASK_D[2][28], ~Iteration_cell_sum_AMASK_D[3][28]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:854:13
				Q_sqrt_com_0 = {{29 {1'b0}}, ~Q_sqrt0[28:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:855:13
				Q_sqrt_com_1 = {{29 {1'b0}}, ~Q_sqrt1[28:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:856:13
				Q_sqrt_com_2 = {{29 {1'b0}}, ~Q_sqrt2[28:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:857:13
				Q_sqrt_com_3 = {{29 {1'b0}}, ~Q_sqrt3[28:0]};
			end
			2'b01: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:861:13
				Sqrt_quotinent_S = {Iteration_cell_carry_D[0], Iteration_cell_carry_D[1], Iteration_cell_carry_D[2], Iteration_cell_carry_D[3]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:862:13
				Q_sqrt_com_0 = ~Q_sqrt0;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:863:13
				Q_sqrt_com_1 = ~Q_sqrt1;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:864:13
				Q_sqrt_com_2 = ~Q_sqrt2;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:865:13
				Q_sqrt_com_3 = ~Q_sqrt3;
			end
			2'b10: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:869:13
				Sqrt_quotinent_S = {~Iteration_cell_sum_AMASK_D[0][15], ~Iteration_cell_sum_AMASK_D[1][15], ~Iteration_cell_sum_AMASK_D[2][15], ~Iteration_cell_sum_AMASK_D[3][15]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:870:13
				Q_sqrt_com_0 = {{42 {1'b0}}, ~Q_sqrt0[15:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:871:13
				Q_sqrt_com_1 = {{42 {1'b0}}, ~Q_sqrt1[15:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:872:13
				Q_sqrt_com_2 = {{42 {1'b0}}, ~Q_sqrt2[15:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:873:13
				Q_sqrt_com_3 = {{42 {1'b0}}, ~Q_sqrt3[15:0]};
			end
			2'b11: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:877:13
				Sqrt_quotinent_S = {~Iteration_cell_sum_AMASK_D[0][12], ~Iteration_cell_sum_AMASK_D[1][12], ~Iteration_cell_sum_AMASK_D[2][12], ~Iteration_cell_sum_AMASK_D[3][12]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:878:13
				Q_sqrt_com_0 = {{45 {1'b0}}, ~Q_sqrt0[12:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:879:13
				Q_sqrt_com_1 = {{45 {1'b0}}, ~Q_sqrt1[12:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:880:13
				Q_sqrt_com_2 = {{45 {1'b0}}, ~Q_sqrt2[12:0]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:881:13
				Q_sqrt_com_3 = {{45 {1'b0}}, ~Q_sqrt3[12:0]};
			end
		endcase
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:888:3
	assign Qcnt_one_0 = 1'b0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:889:3
	assign Qcnt_one_1 = {Quotient_DP[0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:890:3
	assign Qcnt_one_2 = {Quotient_DP[1:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:891:3
	assign Qcnt_one_3 = {Quotient_DP[2:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:892:3
	assign Qcnt_one_4 = {Quotient_DP[3:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:893:3
	assign Qcnt_one_5 = {Quotient_DP[4:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:894:3
	assign Qcnt_one_6 = {Quotient_DP[5:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:895:3
	assign Qcnt_one_7 = {Quotient_DP[6:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:896:3
	assign Qcnt_one_8 = {Quotient_DP[7:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:897:3
	assign Qcnt_one_9 = {Quotient_DP[8:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:898:3
	assign Qcnt_one_10 = {Quotient_DP[9:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:899:3
	assign Qcnt_one_11 = {Quotient_DP[10:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:900:3
	assign Qcnt_one_12 = {Quotient_DP[11:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:901:3
	assign Qcnt_one_13 = {Quotient_DP[12:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:902:3
	assign Qcnt_one_14 = {Quotient_DP[13:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:903:3
	assign Qcnt_one_15 = {Quotient_DP[14:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:904:3
	assign Qcnt_one_16 = {Quotient_DP[15:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:905:3
	assign Qcnt_one_17 = {Quotient_DP[16:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:906:3
	assign Qcnt_one_18 = {Quotient_DP[17:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:907:3
	assign Qcnt_one_19 = {Quotient_DP[18:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:908:3
	assign Qcnt_one_20 = {Quotient_DP[19:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:909:3
	assign Qcnt_one_21 = {Quotient_DP[20:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:910:3
	assign Qcnt_one_22 = {Quotient_DP[21:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:911:3
	assign Qcnt_one_23 = {Quotient_DP[22:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:912:3
	assign Qcnt_one_24 = {Quotient_DP[23:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:913:3
	assign Qcnt_one_25 = {Quotient_DP[24:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:914:3
	assign Qcnt_one_26 = {Quotient_DP[25:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:915:3
	assign Qcnt_one_27 = {Quotient_DP[26:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:916:3
	assign Qcnt_one_28 = {Quotient_DP[27:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:917:3
	assign Qcnt_one_29 = {Quotient_DP[28:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:918:3
	assign Qcnt_one_30 = {Quotient_DP[29:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:919:3
	assign Qcnt_one_31 = {Quotient_DP[30:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:920:3
	assign Qcnt_one_32 = {Quotient_DP[31:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:921:3
	assign Qcnt_one_33 = {Quotient_DP[32:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:922:3
	assign Qcnt_one_34 = {Quotient_DP[33:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:923:3
	assign Qcnt_one_35 = {Quotient_DP[34:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:924:3
	assign Qcnt_one_36 = {Quotient_DP[35:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:925:3
	assign Qcnt_one_37 = {Quotient_DP[36:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:926:3
	assign Qcnt_one_38 = {Quotient_DP[37:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:927:3
	assign Qcnt_one_39 = {Quotient_DP[38:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:928:3
	assign Qcnt_one_40 = {Quotient_DP[39:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:929:3
	assign Qcnt_one_41 = {Quotient_DP[40:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:930:3
	assign Qcnt_one_42 = {Quotient_DP[41:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:931:3
	assign Qcnt_one_43 = {Quotient_DP[42:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:932:3
	assign Qcnt_one_44 = {Quotient_DP[43:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:933:3
	assign Qcnt_one_45 = {Quotient_DP[44:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:934:3
	assign Qcnt_one_46 = {Quotient_DP[45:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:935:3
	assign Qcnt_one_47 = {Quotient_DP[46:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:936:3
	assign Qcnt_one_48 = {Quotient_DP[47:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:937:3
	assign Qcnt_one_49 = {Quotient_DP[48:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:938:3
	assign Qcnt_one_50 = {Quotient_DP[49:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:939:3
	assign Qcnt_one_51 = {Quotient_DP[50:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:940:3
	assign Qcnt_one_52 = {Quotient_DP[51:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:941:3
	assign Qcnt_one_53 = {Quotient_DP[52:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:942:3
	assign Qcnt_one_54 = {Quotient_DP[53:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:943:3
	assign Qcnt_one_55 = {Quotient_DP[54:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:944:3
	assign Qcnt_one_56 = {Quotient_DP[55:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:945:3
	assign Qcnt_one_57 = {Quotient_DP[56:0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:948:3
	assign Qcnt_two_0 = {1'b0, Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:949:3
	assign Qcnt_two_1 = {Quotient_DP[1:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:950:3
	assign Qcnt_two_2 = {Quotient_DP[3:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:951:3
	assign Qcnt_two_3 = {Quotient_DP[5:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:952:3
	assign Qcnt_two_4 = {Quotient_DP[7:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:953:3
	assign Qcnt_two_5 = {Quotient_DP[9:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:954:3
	assign Qcnt_two_6 = {Quotient_DP[11:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:955:3
	assign Qcnt_two_7 = {Quotient_DP[13:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:956:3
	assign Qcnt_two_8 = {Quotient_DP[15:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:957:3
	assign Qcnt_two_9 = {Quotient_DP[17:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:958:3
	assign Qcnt_two_10 = {Quotient_DP[19:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:959:3
	assign Qcnt_two_11 = {Quotient_DP[21:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:960:3
	assign Qcnt_two_12 = {Quotient_DP[23:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:961:3
	assign Qcnt_two_13 = {Quotient_DP[25:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:962:3
	assign Qcnt_two_14 = {Quotient_DP[27:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:963:3
	assign Qcnt_two_15 = {Quotient_DP[29:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:964:3
	assign Qcnt_two_16 = {Quotient_DP[31:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:965:3
	assign Qcnt_two_17 = {Quotient_DP[33:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:966:3
	assign Qcnt_two_18 = {Quotient_DP[35:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:967:3
	assign Qcnt_two_19 = {Quotient_DP[37:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:968:3
	assign Qcnt_two_20 = {Quotient_DP[39:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:969:3
	assign Qcnt_two_21 = {Quotient_DP[41:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:970:3
	assign Qcnt_two_22 = {Quotient_DP[43:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:971:3
	assign Qcnt_two_23 = {Quotient_DP[45:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:972:3
	assign Qcnt_two_24 = {Quotient_DP[47:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:973:3
	assign Qcnt_two_25 = {Quotient_DP[49:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:974:3
	assign Qcnt_two_26 = {Quotient_DP[51:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:975:3
	assign Qcnt_two_27 = {Quotient_DP[53:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:976:3
	assign Qcnt_two_28 = {Quotient_DP[55:0], Sqrt_quotinent_S[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:979:3
	assign Qcnt_three_0 = {1'b0, Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:980:3
	assign Qcnt_three_1 = {Quotient_DP[2:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:981:3
	assign Qcnt_three_2 = {Quotient_DP[5:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:982:3
	assign Qcnt_three_3 = {Quotient_DP[8:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:983:3
	assign Qcnt_three_4 = {Quotient_DP[11:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:984:3
	assign Qcnt_three_5 = {Quotient_DP[14:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:985:3
	assign Qcnt_three_6 = {Quotient_DP[17:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:986:3
	assign Qcnt_three_7 = {Quotient_DP[20:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:987:3
	assign Qcnt_three_8 = {Quotient_DP[23:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:988:3
	assign Qcnt_three_9 = {Quotient_DP[26:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:989:3
	assign Qcnt_three_10 = {Quotient_DP[29:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:990:3
	assign Qcnt_three_11 = {Quotient_DP[32:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:991:3
	assign Qcnt_three_12 = {Quotient_DP[35:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:992:3
	assign Qcnt_three_13 = {Quotient_DP[38:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:993:3
	assign Qcnt_three_14 = {Quotient_DP[41:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:994:3
	assign Qcnt_three_15 = {Quotient_DP[44:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:995:3
	assign Qcnt_three_16 = {Quotient_DP[47:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:996:3
	assign Qcnt_three_17 = {Quotient_DP[50:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:997:3
	assign Qcnt_three_18 = {Quotient_DP[53:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:998:3
	assign Qcnt_three_19 = {Quotient_DP[56:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1001:3
	assign Qcnt_four_0 = {1'b0, Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1002:3
	assign Qcnt_four_1 = {Quotient_DP[3:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1003:3
	assign Qcnt_four_2 = {Quotient_DP[7:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1004:3
	assign Qcnt_four_3 = {Quotient_DP[11:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1005:3
	assign Qcnt_four_4 = {Quotient_DP[15:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1006:3
	assign Qcnt_four_5 = {Quotient_DP[19:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1007:3
	assign Qcnt_four_6 = {Quotient_DP[23:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1008:3
	assign Qcnt_four_7 = {Quotient_DP[27:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1009:3
	assign Qcnt_four_8 = {Quotient_DP[31:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1010:3
	assign Qcnt_four_9 = {Quotient_DP[35:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1011:3
	assign Qcnt_four_10 = {Quotient_DP[39:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1012:3
	assign Qcnt_four_11 = {Quotient_DP[43:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1013:3
	assign Qcnt_four_12 = {Quotient_DP[47:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1014:3
	assign Qcnt_four_13 = {Quotient_DP[51:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1015:3
	assign Qcnt_four_14 = {Quotient_DP[55:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1020:3
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1022:3
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1033:9
				case (Crtl_cnt_S)
					6'b000000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1037:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1038:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_one_0};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1039:15
						Sqrt_Q0 = Q_sqrt_com_0;
					end
					6'b000001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1043:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[51:50];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1044:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_one_1};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1045:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1049:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[49:48];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1050:15
						Q_sqrt0 = {{56 {1'b0}}, Qcnt_one_2};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1051:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1055:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[47:46];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1056:15
						Q_sqrt0 = {{55 {1'b0}}, Qcnt_one_3};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1057:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1061:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[45:44];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1062:15
						Q_sqrt0 = {{54 {1'b0}}, Qcnt_one_4};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1063:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1067:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[43:42];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1068:15
						Q_sqrt0 = {{53 {1'b0}}, Qcnt_one_5};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1069:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1073:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[41:40];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1074:15
						Q_sqrt0 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_one_6};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1075:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1079:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[39:38];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1080:15
						Q_sqrt0 = {{51 {1'b0}}, Qcnt_one_7};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1081:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1085:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[37:36];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1086:15
						Q_sqrt0 = {{50 {1'b0}}, Qcnt_one_8};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1087:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1091:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[35:34];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1092:15
						Q_sqrt0 = {{49 {1'b0}}, Qcnt_one_9};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1093:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1097:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[33:32];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1098:15
						Q_sqrt0 = {{48 {1'b0}}, Qcnt_one_10};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1099:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1103:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[31:30];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1104:15
						Q_sqrt0 = {{47 {1'b0}}, Qcnt_one_11};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1105:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1109:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1110:15
						Q_sqrt0 = {{46 {1'b0}}, Qcnt_one_12};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1111:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1115:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[27:26];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1116:15
						Q_sqrt0 = {{45 {1'b0}}, Qcnt_one_13};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1117:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1121:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[25:24];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1122:15
						Q_sqrt0 = {{44 {1'b0}}, Qcnt_one_14};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1123:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1127:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[23:22];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1128:15
						Q_sqrt0 = {{43 {1'b0}}, Qcnt_one_15};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1129:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1133:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[21:20];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1134:15
						Q_sqrt0 = {{42 {1'b0}}, Qcnt_one_16};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1135:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1139:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[19:18];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1140:15
						Q_sqrt0 = {{41 {1'b0}}, Qcnt_one_17};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1141:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1145:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[17:16];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1146:15
						Q_sqrt0 = {{40 {1'b0}}, Qcnt_one_18};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1147:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1151:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[15:14];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1152:15
						Q_sqrt0 = {{39 {1'b0}}, Qcnt_one_19};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1153:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1157:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[13:12];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1158:15
						Q_sqrt0 = {{38 {1'b0}}, Qcnt_one_20};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1159:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1163:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[11:10];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1164:15
						Q_sqrt0 = {{37 {1'b0}}, Qcnt_one_21};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1165:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1169:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[9:8];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1170:15
						Q_sqrt0 = {{36 {1'b0}}, Qcnt_one_22};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1171:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1175:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[7:6];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1176:15
						Q_sqrt0 = {{35 {1'b0}}, Qcnt_one_23};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1177:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1181:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1182:15
						Q_sqrt0 = {{34 {1'b0}}, Qcnt_one_24};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1183:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1187:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[3:2];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1188:15
						Q_sqrt0 = {{33 {1'b0}}, Qcnt_one_25};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1189:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1193:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[1:0];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1194:15
						Q_sqrt0 = {{32 {1'b0}}, Qcnt_one_26};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1195:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1199:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1200:15
						Q_sqrt0 = {{31 {1'b0}}, Qcnt_one_27};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1201:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1205:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1206:15
						Q_sqrt0 = {{30 {1'b0}}, Qcnt_one_28};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1207:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1211:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1212:15
						Q_sqrt0 = {{29 {1'b0}}, Qcnt_one_29};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1213:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1217:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1218:15
						Q_sqrt0 = {{28 {1'b0}}, Qcnt_one_30};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1219:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1223:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1224:15
						Q_sqrt0 = {{27 {1'b0}}, Qcnt_one_31};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1225:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1229:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1230:15
						Q_sqrt0 = {{26 {1'b0}}, Qcnt_one_32};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1231:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1235:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1236:15
						Q_sqrt0 = {{25 {1'b0}}, Qcnt_one_33};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1237:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1241:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1242:15
						Q_sqrt0 = {{24 {1'b0}}, Qcnt_one_34};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1243:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1247:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1248:15
						Q_sqrt0 = {{23 {1'b0}}, Qcnt_one_35};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1249:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1253:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1254:15
						Q_sqrt0 = {{22 {1'b0}}, Qcnt_one_36};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1255:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1259:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1260:15
						Q_sqrt0 = {{21 {1'b0}}, Qcnt_one_37};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1261:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1265:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1266:15
						Q_sqrt0 = {{20 {1'b0}}, Qcnt_one_38};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1267:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1271:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1272:15
						Q_sqrt0 = {{19 {1'b0}}, Qcnt_one_39};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1273:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1277:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1278:15
						Q_sqrt0 = {{18 {1'b0}}, Qcnt_one_40};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1279:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1283:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1284:15
						Q_sqrt0 = {{17 {1'b0}}, Qcnt_one_41};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1285:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1289:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1290:15
						Q_sqrt0 = {{16 {1'b0}}, Qcnt_one_42};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1291:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1295:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1296:15
						Q_sqrt0 = {{15 {1'b0}}, Qcnt_one_43};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1297:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1301:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1302:15
						Q_sqrt0 = {{14 {1'b0}}, Qcnt_one_44};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1303:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1307:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1308:15
						Q_sqrt0 = {{13 {1'b0}}, Qcnt_one_45};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1309:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1313:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1314:15
						Q_sqrt0 = {{12 {1'b0}}, Qcnt_one_46};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1315:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1319:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1320:15
						Q_sqrt0 = {{11 {1'b0}}, Qcnt_one_47};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1321:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1325:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1326:15
						Q_sqrt0 = {{10 {1'b0}}, Qcnt_one_48};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1327:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1331:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1332:15
						Q_sqrt0 = {{9 {1'b0}}, Qcnt_one_49};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1333:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1337:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1338:15
						Q_sqrt0 = {{8 {1'b0}}, Qcnt_one_50};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1339:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1343:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1344:15
						Q_sqrt0 = {{7 {1'b0}}, Qcnt_one_51};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1345:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1349:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1350:15
						Q_sqrt0 = {{6 {1'b0}}, Qcnt_one_52};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1351:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1355:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1356:15
						Q_sqrt0 = {{5 {1'b0}}, Qcnt_one_53};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1357:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1361:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1362:15
						Q_sqrt0 = {{4 {1'b0}}, Qcnt_one_54};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1363:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1367:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1368:15
						Q_sqrt0 = {{3 {1'b0}}, Qcnt_one_55};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1369:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b111000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1373:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1374:15
						Q_sqrt0 = {{2 {1'b0}}, Qcnt_one_56};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1375:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					default: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1380:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1381:15
						Q_sqrt0 = 1'sb0;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1382:15
						Sqrt_Q0 = 1'sb0;
					end
				endcase
			2'b01:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1398:9
				case (Crtl_cnt_S)
					6'b000000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1402:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1403:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_two_0[1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1404:15
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1405:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1406:15
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_two_0[1:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1407:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1412:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[49:48];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1413:15
						Q_sqrt0 = {{56 {1'b0}}, Qcnt_two_1[2:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1414:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1415:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[47:46];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1416:15
						Q_sqrt1 = {{55 {1'b0}}, Qcnt_two_1[2:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1417:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1422:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[45:44];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1423:15
						Q_sqrt0 = {{54 {1'b0}}, Qcnt_two_2[4:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1424:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1425:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[43:42];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1426:15
						Q_sqrt1 = {{53 {1'b0}}, Qcnt_two_2[4:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1427:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1432:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[41:40];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1433:15
						Q_sqrt0 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_two_3[6:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1434:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1435:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[39:38];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1436:15
						Q_sqrt1 = {{51 {1'b0}}, Qcnt_two_3[6:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1437:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1442:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[37:36];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1443:15
						Q_sqrt0 = {{50 {1'b0}}, Qcnt_two_4[8:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1444:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1445:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[35:34];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1446:15
						Q_sqrt1 = {{49 {1'b0}}, Qcnt_two_4[8:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1447:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1452:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[33:32];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1453:15
						Q_sqrt0 = {{48 {1'b0}}, Qcnt_two_5[10:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1454:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1455:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[31:30];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1456:15
						Q_sqrt1 = {{47 {1'b0}}, Qcnt_two_5[10:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1457:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1462:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1463:15
						Q_sqrt0 = {{46 {1'b0}}, Qcnt_two_6[12:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1464:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1465:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[27:26];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1466:15
						Q_sqrt1 = {{45 {1'b0}}, Qcnt_two_6[12:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1467:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1472:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[25:24];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1473:15
						Q_sqrt0 = {{44 {1'b0}}, Qcnt_two_7[14:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1474:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1475:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[23:22];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1476:15
						Q_sqrt1 = {{43 {1'b0}}, Qcnt_two_7[14:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1477:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1482:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[21:20];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1483:15
						Q_sqrt0 = {{42 {1'b0}}, Qcnt_two_8[16:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1484:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1485:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[19:18];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1486:15
						Q_sqrt1 = {{41 {1'b0}}, Qcnt_two_8[16:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1487:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1492:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[17:16];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1493:15
						Q_sqrt0 = {{40 {1'b0}}, Qcnt_two_9[18:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1494:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1495:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[15:14];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1496:15
						Q_sqrt1 = {{39 {1'b0}}, Qcnt_two_9[18:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1497:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1502:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[13:12];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1503:15
						Q_sqrt0 = {{38 {1'b0}}, Qcnt_two_10[20:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1504:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1505:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[11:10];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1506:15
						Q_sqrt1 = {{37 {1'b0}}, Qcnt_two_10[20:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1507:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1512:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[9:8];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1513:15
						Q_sqrt0 = {{36 {1'b0}}, Qcnt_two_11[22:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1514:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1515:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[7:6];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1516:15
						Q_sqrt1 = {{35 {1'b0}}, Qcnt_two_11[22:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1517:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1522:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1523:15
						Q_sqrt0 = {{34 {1'b0}}, Qcnt_two_12[24:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1524:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1525:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[3:2];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1526:15
						Q_sqrt1 = {{33 {1'b0}}, Qcnt_two_12[24:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1527:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1532:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[1:0];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1533:15
						Q_sqrt0 = {{32 {1'b0}}, Qcnt_two_13[26:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1534:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1535:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1536:15
						Q_sqrt1 = {{31 {1'b0}}, Qcnt_two_13[26:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1537:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1542:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1543:15
						Q_sqrt0 = {{30 {1'b0}}, Qcnt_two_14[28:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1544:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1545:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1546:15
						Q_sqrt1 = {{29 {1'b0}}, Qcnt_two_14[28:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1547:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1552:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1553:15
						Q_sqrt0 = {{28 {1'b0}}, Qcnt_two_15[30:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1554:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1555:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1556:15
						Q_sqrt1 = {{27 {1'b0}}, Qcnt_two_15[30:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1557:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1562:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1563:15
						Q_sqrt0 = {{26 {1'b0}}, Qcnt_two_16[32:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1564:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1565:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1566:15
						Q_sqrt1 = {{25 {1'b0}}, Qcnt_two_16[32:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1567:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1572:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1573:15
						Q_sqrt0 = {{24 {1'b0}}, Qcnt_two_17[34:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1574:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1575:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1576:15
						Q_sqrt1 = {{23 {1'b0}}, Qcnt_two_17[34:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1577:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1582:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1583:15
						Q_sqrt0 = {{22 {1'b0}}, Qcnt_two_18[36:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1584:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1585:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1586:15
						Q_sqrt1 = {{21 {1'b0}}, Qcnt_two_18[36:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1587:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1592:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1593:15
						Q_sqrt0 = {{20 {1'b0}}, Qcnt_two_19[38:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1594:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1595:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1596:15
						Q_sqrt1 = {{19 {1'b0}}, Qcnt_two_19[38:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1597:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1602:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1603:15
						Q_sqrt0 = {{18 {1'b0}}, Qcnt_two_20[40:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1604:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1605:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1606:15
						Q_sqrt1 = {{17 {1'b0}}, Qcnt_two_20[40:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1607:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1612:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1613:15
						Q_sqrt0 = {{16 {1'b0}}, Qcnt_two_21[42:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1614:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1615:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1616:15
						Q_sqrt1 = {{15 {1'b0}}, Qcnt_two_21[42:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1617:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1622:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1623:15
						Q_sqrt0 = {{14 {1'b0}}, Qcnt_two_22[44:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1624:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1625:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1626:15
						Q_sqrt1 = {{13 {1'b0}}, Qcnt_two_22[44:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1627:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1632:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1633:15
						Q_sqrt0 = {{12 {1'b0}}, Qcnt_two_23[46:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1634:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1635:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1636:15
						Q_sqrt1 = {{11 {1'b0}}, Qcnt_two_23[46:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1637:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1642:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1643:15
						Q_sqrt0 = {{10 {1'b0}}, Qcnt_two_24[48:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1644:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1645:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1646:15
						Q_sqrt1 = {{9 {1'b0}}, Qcnt_two_24[48:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1647:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1652:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1653:15
						Q_sqrt0 = {{8 {1'b0}}, Qcnt_two_25[50:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1654:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1655:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1656:15
						Q_sqrt1 = {{7 {1'b0}}, Qcnt_two_25[50:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1657:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1662:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1663:15
						Q_sqrt0 = {{6 {1'b0}}, Qcnt_two_26[52:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1664:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1665:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1666:15
						Q_sqrt1 = {{5 {1'b0}}, Qcnt_two_26[52:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1667:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1672:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1673:15
						Q_sqrt0 = {{4 {1'b0}}, Qcnt_two_27[54:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1674:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1675:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1676:15
						Q_sqrt1 = {{3 {1'b0}}, Qcnt_two_27[54:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1677:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1682:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1683:15
						Q_sqrt0 = {{2 {1'b0}}, Qcnt_two_28[56:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1684:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1685:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1686:15
						Q_sqrt1 = {1'b0, Qcnt_two_28[56:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1687:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					default: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1692:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1693:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_two_0[1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1694:15
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1695:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1696:15
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_two_0[1:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1697:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
				endcase
			2'b10:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1714:9
				case (Crtl_cnt_S)
					6'b000000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1717:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1718:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_three_0[2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1719:15
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1720:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1721:15
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_three_0[2:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1722:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1723:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1724:15
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_three_0[2:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1725:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1730:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[47:46];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1731:15
						Q_sqrt0 = {{54 {1'b0}}, Qcnt_three_1[4:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1732:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1733:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[45:44];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1734:15
						Q_sqrt1 = {{53 {1'b0}}, Qcnt_three_1[4:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1735:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1736:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[43:42];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1737:15
						Q_sqrt2 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_three_1[4:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1738:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1743:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[41:40];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1744:15
						Q_sqrt0 = {{51 {1'b0}}, Qcnt_three_2[7:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1745:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1746:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[39:38];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1747:15
						Q_sqrt1 = {{50 {1'b0}}, Qcnt_three_2[7:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1748:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1749:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[37:36];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1750:15
						Q_sqrt2 = {{49 {1'b0}}, Qcnt_three_2[7:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1751:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1756:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[35:34];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1757:15
						Q_sqrt0 = {{48 {1'b0}}, Qcnt_three_3[10:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1758:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1759:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[33:32];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1760:15
						Q_sqrt1 = {{47 {1'b0}}, Qcnt_three_3[10:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1761:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1762:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[31:30];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1763:15
						Q_sqrt2 = {{46 {1'b0}}, Qcnt_three_3[10:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1764:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1769:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1770:15
						Q_sqrt0 = {{45 {1'b0}}, Qcnt_three_4[13:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1771:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1772:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[27:26];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1773:15
						Q_sqrt1 = {{44 {1'b0}}, Qcnt_three_4[13:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1774:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1775:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[25:24];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1776:15
						Q_sqrt2 = {{43 {1'b0}}, Qcnt_three_4[13:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1777:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1782:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[23:22];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1783:15
						Q_sqrt0 = {{42 {1'b0}}, Qcnt_three_5[16:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1784:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1785:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[21:20];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1786:15
						Q_sqrt1 = {{41 {1'b0}}, Qcnt_three_5[16:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1787:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1788:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[19:18];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1789:15
						Q_sqrt2 = {{40 {1'b0}}, Qcnt_three_5[16:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1790:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1795:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[17:16];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1796:15
						Q_sqrt0 = {{39 {1'b0}}, Qcnt_three_6[19:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1797:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1798:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[15:14];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1799:15
						Q_sqrt1 = {{38 {1'b0}}, Qcnt_three_6[19:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1800:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1801:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[13:12];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1802:15
						Q_sqrt2 = {{37 {1'b0}}, Qcnt_three_6[19:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1803:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1808:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[11:10];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1809:15
						Q_sqrt0 = {{36 {1'b0}}, Qcnt_three_7[22:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1810:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1811:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[9:8];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1812:15
						Q_sqrt1 = {{35 {1'b0}}, Qcnt_three_7[22:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1813:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1814:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[7:6];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1815:15
						Q_sqrt2 = {{34 {1'b0}}, Qcnt_three_7[22:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1816:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1821:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1822:15
						Q_sqrt0 = {{33 {1'b0}}, Qcnt_three_8[25:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1823:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1824:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[3:2];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1825:15
						Q_sqrt1 = {{32 {1'b0}}, Qcnt_three_8[25:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1826:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1827:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[1:0];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1828:15
						Q_sqrt2 = {{31 {1'b0}}, Qcnt_three_8[25:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1829:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1834:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1835:15
						Q_sqrt0 = {{30 {1'b0}}, Qcnt_three_9[28:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1836:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1837:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1838:15
						Q_sqrt1 = {{29 {1'b0}}, Qcnt_three_9[28:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1839:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1840:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1841:15
						Q_sqrt2 = {{28 {1'b0}}, Qcnt_three_9[28:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1842:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1847:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1848:15
						Q_sqrt0 = {{27 {1'b0}}, Qcnt_three_10[31:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1849:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1850:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1851:15
						Q_sqrt1 = {{26 {1'b0}}, Qcnt_three_10[31:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1852:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1853:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1854:15
						Q_sqrt2 = {{25 {1'b0}}, Qcnt_three_10[31:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1855:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1860:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1861:15
						Q_sqrt0 = {{24 {1'b0}}, Qcnt_three_11[34:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1862:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1863:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1864:15
						Q_sqrt1 = {{23 {1'b0}}, Qcnt_three_11[34:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1865:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1866:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1867:15
						Q_sqrt2 = {{22 {1'b0}}, Qcnt_three_11[34:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1868:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1873:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1874:15
						Q_sqrt0 = {{21 {1'b0}}, Qcnt_three_12[37:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1875:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1876:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1877:15
						Q_sqrt1 = {{20 {1'b0}}, Qcnt_three_12[37:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1878:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1879:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1880:15
						Q_sqrt2 = {{19 {1'b0}}, Qcnt_three_12[37:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1881:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1886:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1887:15
						Q_sqrt0 = {{18 {1'b0}}, Qcnt_three_13[40:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1888:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1889:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1890:15
						Q_sqrt1 = {{17 {1'b0}}, Qcnt_three_13[40:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1891:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1892:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1893:15
						Q_sqrt2 = {{16 {1'b0}}, Qcnt_three_13[40:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1894:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1899:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1900:15
						Q_sqrt0 = {{15 {1'b0}}, Qcnt_three_14[43:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1901:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1902:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1903:15
						Q_sqrt1 = {{14 {1'b0}}, Qcnt_three_14[43:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1904:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1905:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1906:15
						Q_sqrt2 = {{13 {1'b0}}, Qcnt_three_14[43:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1907:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1912:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1913:15
						Q_sqrt0 = {{12 {1'b0}}, Qcnt_three_15[46:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1914:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1915:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1916:15
						Q_sqrt1 = {{11 {1'b0}}, Qcnt_three_15[46:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1917:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1918:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1919:15
						Q_sqrt2 = {{10 {1'b0}}, Qcnt_three_15[46:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1920:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b010000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1925:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1926:15
						Q_sqrt0 = {{9 {1'b0}}, Qcnt_three_16[49:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1927:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1928:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1929:15
						Q_sqrt1 = {{8 {1'b0}}, Qcnt_three_16[49:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1930:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1931:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1932:15
						Q_sqrt2 = {{7 {1'b0}}, Qcnt_three_16[49:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1933:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b010001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1938:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1939:15
						Q_sqrt0 = {{6 {1'b0}}, Qcnt_three_17[52:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1940:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1941:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1942:15
						Q_sqrt1 = {{5 {1'b0}}, Qcnt_three_17[52:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1943:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1944:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1945:15
						Q_sqrt2 = {{4 {1'b0}}, Qcnt_three_17[52:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1946:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b010010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1951:15
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1952:15
						Q_sqrt0 = {{3 {1'b0}}, Qcnt_three_18[55:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1953:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1954:15
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1955:15
						Q_sqrt1 = {{2 {1'b0}}, Qcnt_three_18[55:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1956:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1957:15
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1958:15
						Q_sqrt2 = {1'b0, Qcnt_three_18[55:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1959:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					default: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1964:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1965:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_three_0[2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1966:15
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1967:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1968:15
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_three_0[2:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1969:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1970:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1971:15
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_three_0[2:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1972:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
				endcase
			2'b11:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1988:15
				case (Crtl_cnt_S)
					6'b000000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1992:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1993:21
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_four_0[3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1994:21
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1995:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1996:21
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_four_0[3:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1997:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1998:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1999:21
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_four_0[3:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2000:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2001:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[47:46];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2002:21
						Q_sqrt3 = {{54 {1'b0}}, Qcnt_four_0[3:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2003:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2008:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[45:44];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2009:21
						Q_sqrt0 = {{53 {1'b0}}, Qcnt_four_1[6:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2010:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2011:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[43:42];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2012:21
						Q_sqrt1 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_four_1[6:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2013:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2014:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[41:40];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2015:21
						Q_sqrt2 = {{51 {1'b0}}, Qcnt_four_1[6:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2016:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2017:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[39:38];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2018:21
						Q_sqrt3 = {{50 {1'b0}}, Qcnt_four_1[6:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2019:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2024:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[37:36];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2025:21
						Q_sqrt0 = {{49 {1'b0}}, Qcnt_four_2[10:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2026:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2027:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[35:34];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2028:21
						Q_sqrt1 = {{48 {1'b0}}, Qcnt_four_2[10:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2029:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2030:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[33:32];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2031:21
						Q_sqrt2 = {{47 {1'b0}}, Qcnt_four_2[10:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2032:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2033:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[31:30];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2034:21
						Q_sqrt3 = {{46 {1'b0}}, Qcnt_four_2[10:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2035:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2040:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2041:21
						Q_sqrt0 = {{45 {1'b0}}, Qcnt_four_3[14:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2042:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2043:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[27:26];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2044:21
						Q_sqrt1 = {{44 {1'b0}}, Qcnt_four_3[14:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2045:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2046:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[25:24];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2047:21
						Q_sqrt2 = {{43 {1'b0}}, Qcnt_four_3[14:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2048:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2049:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[23:22];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2050:21
						Q_sqrt3 = {{42 {1'b0}}, Qcnt_four_3[14:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2051:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2056:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[21:20];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2057:21
						Q_sqrt0 = {{41 {1'b0}}, Qcnt_four_4[18:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2058:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2059:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[19:18];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2060:21
						Q_sqrt1 = {{40 {1'b0}}, Qcnt_four_4[18:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2061:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2062:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[17:16];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2063:21
						Q_sqrt2 = {{39 {1'b0}}, Qcnt_four_4[18:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2064:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2065:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[15:14];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2066:21
						Q_sqrt3 = {{38 {1'b0}}, Qcnt_four_4[18:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2067:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2072:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[13:12];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2073:21
						Q_sqrt0 = {{37 {1'b0}}, Qcnt_four_5[22:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2074:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2075:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[11:10];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2076:21
						Q_sqrt1 = {{36 {1'b0}}, Qcnt_four_5[22:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2077:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2078:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[9:8];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2079:21
						Q_sqrt2 = {{35 {1'b0}}, Qcnt_four_5[22:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2080:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2081:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[7:6];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2082:21
						Q_sqrt3 = {{34 {1'b0}}, Qcnt_four_5[22:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2083:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000110: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2088:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2089:21
						Q_sqrt0 = {{33 {1'b0}}, Qcnt_four_6[26:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2090:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2091:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[3:2];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2092:21
						Q_sqrt1 = {{32 {1'b0}}, Qcnt_four_6[26:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2093:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2094:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[1:0];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2095:21
						Q_sqrt2 = {{31 {1'b0}}, Qcnt_four_6[26:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2096:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2097:21
						Sqrt_DI[3] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2098:21
						Q_sqrt3 = {{30 {1'b0}}, Qcnt_four_6[26:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2099:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000111: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2104:21
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2105:21
						Q_sqrt0 = {{29 {1'b0}}, Qcnt_four_7[30:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2106:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2107:21
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2108:21
						Q_sqrt1 = {{28 {1'b0}}, Qcnt_four_7[30:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2109:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2110:21
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2111:21
						Q_sqrt2 = {{27 {1'b0}}, Qcnt_four_7[30:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2112:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2113:21
						Sqrt_DI[3] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2114:21
						Q_sqrt3 = {{26 {1'b0}}, Qcnt_four_7[30:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2115:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001000: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2120:21
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2121:21
						Q_sqrt0 = {{25 {1'b0}}, Qcnt_four_8[34:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2122:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2123:21
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2124:21
						Q_sqrt1 = {{24 {1'b0}}, Qcnt_four_8[34:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2125:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2126:21
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2127:21
						Q_sqrt2 = {{23 {1'b0}}, Qcnt_four_8[34:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2128:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2129:21
						Sqrt_DI[3] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2130:21
						Q_sqrt3 = {{22 {1'b0}}, Qcnt_four_8[34:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2131:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001001: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2136:21
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2137:21
						Q_sqrt0 = {{21 {1'b0}}, Qcnt_four_9[38:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2138:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2139:21
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2140:21
						Q_sqrt1 = {{20 {1'b0}}, Qcnt_four_9[38:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2141:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2142:21
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2143:21
						Q_sqrt2 = {{19 {1'b0}}, Qcnt_four_9[38:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2144:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2145:21
						Sqrt_DI[3] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2146:21
						Q_sqrt3 = {{18 {1'b0}}, Qcnt_four_9[38:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2147:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001010: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2152:21
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2153:21
						Q_sqrt0 = {{17 {1'b0}}, Qcnt_four_10[42:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2154:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2155:21
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2156:21
						Q_sqrt1 = {{16 {1'b0}}, Qcnt_four_10[42:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2157:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2158:21
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2159:21
						Q_sqrt2 = {{15 {1'b0}}, Qcnt_four_10[42:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2160:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2161:21
						Sqrt_DI[3] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2162:21
						Q_sqrt3 = {{14 {1'b0}}, Qcnt_four_10[42:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2163:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001011: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2168:21
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2169:21
						Q_sqrt0 = {{13 {1'b0}}, Qcnt_four_11[46:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2170:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2171:21
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2172:21
						Q_sqrt1 = {{12 {1'b0}}, Qcnt_four_11[46:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2173:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2174:21
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2175:21
						Q_sqrt2 = {{11 {1'b0}}, Qcnt_four_11[46:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2176:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2177:21
						Sqrt_DI[3] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2178:21
						Q_sqrt3 = {{10 {1'b0}}, Qcnt_four_11[46:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2179:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001100: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2184:21
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2185:21
						Q_sqrt0 = {{9 {1'b0}}, Qcnt_four_12[50:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2186:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2187:21
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2188:21
						Q_sqrt1 = {{8 {1'b0}}, Qcnt_four_12[50:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2189:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2190:21
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2191:21
						Q_sqrt2 = {{7 {1'b0}}, Qcnt_four_12[50:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2192:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2193:21
						Sqrt_DI[3] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2194:21
						Q_sqrt3 = {{6 {1'b0}}, Qcnt_four_12[50:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2195:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001101: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2200:21
						Sqrt_DI[0] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2201:21
						Q_sqrt0 = {{5 {1'b0}}, Qcnt_four_13[54:3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2202:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2203:21
						Sqrt_DI[1] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2204:21
						Q_sqrt1 = {{4 {1'b0}}, Qcnt_four_13[54:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2205:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2206:21
						Sqrt_DI[2] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2207:21
						Q_sqrt2 = {{3 {1'b0}}, Qcnt_four_13[54:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2208:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2209:21
						Sqrt_DI[3] = 2'b00;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2210:21
						Q_sqrt3 = {{2 {1'b0}}, Qcnt_four_13[54:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2211:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					default: begin
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2216:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2217:21
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_four_0[3]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2218:21
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2219:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2220:21
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_four_0[3:2]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2221:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2222:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2223:21
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_four_0[3:1]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2224:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2225:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[47:46];
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2226:21
						Q_sqrt3 = {{54 {1'b0}}, Qcnt_four_0[3:0]};
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2227:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
				endcase
		endcase
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2239:3
	assign Sqrt_R0 = (Sqrt_start_dly_S ? {58 {1'sb0}} : {Partial_remainder_DP[57:0]});
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2240:3
	assign Sqrt_R1 = {Iteration_cell_sum_AMASK_D[0][57], Iteration_cell_sum_AMASK_D[0][54:0], Sqrt_DO[0]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2241:3
	assign Sqrt_R2 = {Iteration_cell_sum_AMASK_D[1][57], Iteration_cell_sum_AMASK_D[1][54:0], Sqrt_DO[1]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2242:3
	assign Sqrt_R3 = {Iteration_cell_sum_AMASK_D[2][57], Iteration_cell_sum_AMASK_D[2][54:0], Sqrt_DO[2]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2243:3
	assign Sqrt_R4 = {Iteration_cell_sum_AMASK_D[3][57], Iteration_cell_sum_AMASK_D[3][54:0], Sqrt_DO[3]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2245:3
	wire [57:0] Denominator_se_format_DB;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2247:3
	assign Denominator_se_format_DB = {Denominator_se_DB[53:45], (FP16ALT_SO ? FP16ALT_SO : Denominator_se_DB[44]), Denominator_se_DB[43:42], (FP16_SO ? FP16_SO : Denominator_se_DB[41]), Denominator_se_DB[40:29], (FP32_SO ? FP32_SO : Denominator_se_DB[28]), Denominator_se_DB[27:0], FP64_SO, 3'b000};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2252:3
	wire [57:0] First_iteration_cell_div_a_D;
	wire [57:0] First_iteration_cell_div_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2253:3
	wire Sel_b_for_first_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2256:3
	assign First_iteration_cell_div_a_D = (Div_start_dly_S ? {Numerator_se_D[53:45], (FP16ALT_SO ? FP16ALT_SO : Numerator_se_D[44]), Numerator_se_D[43:42], (FP16_SO ? FP16_SO : Numerator_se_D[41]), Numerator_se_D[40:29], (FP32_SO ? FP32_SO : Numerator_se_D[28]), Numerator_se_D[27:0], FP64_SO, 3'b000} : {Partial_remainder_DP[56:48], (FP16ALT_SO ? Quotient_DP[0] : Partial_remainder_DP[47]), Partial_remainder_DP[46:45], (FP16_SO ? Quotient_DP[0] : Partial_remainder_DP[44]), Partial_remainder_DP[43:32], (FP32_SO ? Quotient_DP[0] : Partial_remainder_DP[31]), Partial_remainder_DP[30:3], FP64_SO && Quotient_DP[0], 3'b000});
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2264:3
	assign Sel_b_for_first_S = (Div_start_dly_S ? 1 : Quotient_DP[0]);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2265:3
	assign First_iteration_cell_div_b_D = (Sel_b_for_first_S ? Denominator_se_format_DB : {Denominator_se_D, 4'b0000});
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2266:3
	assign Iteration_cell_a_BMASK_D[0] = (Sqrt_enable_SO ? Sqrt_R0 : {First_iteration_cell_div_a_D});
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2267:3
	assign Iteration_cell_b_BMASK_D[0] = (Sqrt_enable_SO ? Sqrt_Q0 : {First_iteration_cell_div_b_D});
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2272:3
	wire [57:0] Sec_iteration_cell_div_a_D;
	wire [57:0] Sec_iteration_cell_div_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2273:3
	wire Sel_b_for_sec_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2274:3
	generate
		if (|defs_div_sqrt_mvp_Iteration_unit_num_S) begin : genblk1
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2277:9
			assign Sel_b_for_sec_S = ~Iteration_cell_sum_AMASK_D[0][57];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2278:9
			assign Sec_iteration_cell_div_a_D = {Iteration_cell_sum_AMASK_D[0][56:48], (FP16ALT_SO ? Sel_b_for_sec_S : Iteration_cell_sum_AMASK_D[0][47]), Iteration_cell_sum_AMASK_D[0][46:45], (FP16_SO ? Sel_b_for_sec_S : Iteration_cell_sum_AMASK_D[0][44]), Iteration_cell_sum_AMASK_D[0][43:32], (FP32_SO ? Sel_b_for_sec_S : Iteration_cell_sum_AMASK_D[0][31]), Iteration_cell_sum_AMASK_D[0][30:3], FP64_SO && Sel_b_for_sec_S, 3'b000};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2282:9
			assign Sec_iteration_cell_div_b_D = (Sel_b_for_sec_S ? Denominator_se_format_DB : {Denominator_se_D, 4'b0000});
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2283:9
			assign Iteration_cell_a_BMASK_D[1] = (Sqrt_enable_SO ? Sqrt_R1 : {Sec_iteration_cell_div_a_D});
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2284:9
			assign Iteration_cell_b_BMASK_D[1] = (Sqrt_enable_SO ? Sqrt_Q1 : {Sec_iteration_cell_div_b_D});
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2289:3
	wire [57:0] Thi_iteration_cell_div_a_D;
	wire [57:0] Thi_iteration_cell_div_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2290:3
	wire Sel_b_for_thi_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2291:3
	generate
		if (1'd1 | 1'd0) begin : genblk2
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2294:9
			assign Sel_b_for_thi_S = ~Iteration_cell_sum_AMASK_D[1][57];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2295:9
			assign Thi_iteration_cell_div_a_D = {Iteration_cell_sum_AMASK_D[1][56:48], (FP16ALT_SO ? Sel_b_for_thi_S : Iteration_cell_sum_AMASK_D[1][47]), Iteration_cell_sum_AMASK_D[1][46:45], (FP16_SO ? Sel_b_for_thi_S : Iteration_cell_sum_AMASK_D[1][44]), Iteration_cell_sum_AMASK_D[1][43:32], (FP32_SO ? Sel_b_for_thi_S : Iteration_cell_sum_AMASK_D[1][31]), Iteration_cell_sum_AMASK_D[1][30:3], FP64_SO && Sel_b_for_thi_S, 3'b000};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2299:9
			assign Thi_iteration_cell_div_b_D = (Sel_b_for_thi_S ? Denominator_se_format_DB : {Denominator_se_D, 4'b0000});
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2300:9
			assign Iteration_cell_a_BMASK_D[2] = (Sqrt_enable_SO ? Sqrt_R2 : {Thi_iteration_cell_div_a_D});
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2301:9
			assign Iteration_cell_b_BMASK_D[2] = (Sqrt_enable_SO ? Sqrt_Q2 : {Thi_iteration_cell_div_b_D});
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2306:3
	wire [57:0] Fou_iteration_cell_div_a_D;
	wire [57:0] Fou_iteration_cell_div_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2307:3
	wire Sel_b_for_fou_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2309:3
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2328:3
	wire [57:0] Mask_bits_ctl_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2330:3
	assign Mask_bits_ctl_S = 58'h3ffffffffffffff;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2337:3
	wire Div_enable_SI [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2338:3
	wire Div_start_dly_SI [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2339:3
	wire Sqrt_enable_SI [3:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2340:3
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2341:5
	genvar _gv_i_265;
	genvar _gv_j_30;
	generate
		for (_gv_i_265 = 0; _gv_i_265 <= defs_div_sqrt_mvp_Iteration_unit_num_S; _gv_i_265 = _gv_i_265 + 1) begin : genblk4
			localparam i = _gv_i_265;
			for (_gv_j_30 = 0; _gv_j_30 <= 57; _gv_j_30 = _gv_j_30 + 1) begin : genblk1
				localparam j = _gv_j_30;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2345:15
				assign Iteration_cell_a_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_a_BMASK_D[i][j];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2346:15
				assign Iteration_cell_b_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_b_BMASK_D[i][j];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2347:15
				assign Iteration_cell_sum_AMASK_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_sum_D[i][j];
			end
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2350:11
			assign Div_enable_SI[i] = Div_enable_SO;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2351:11
			assign Div_start_dly_SI[i] = Div_start_dly_S;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2352:11
			assign Sqrt_enable_SI[i] = Sqrt_enable_SO;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2353:11
			iteration_div_sqrt_mvp #(.WIDTH(58)) iteration_div_sqrt(
				.A_DI(Iteration_cell_a_D[i]),
				.B_DI(Iteration_cell_b_D[i]),
				.Div_enable_SI(Div_enable_SI[i]),
				.Div_start_dly_SI(Div_start_dly_SI[i]),
				.Sqrt_enable_SI(Sqrt_enable_SI[i]),
				.D_DI(Sqrt_DI[i]),
				.D_DO(Sqrt_DO[i]),
				.Sum_DO(Iteration_cell_sum_D[i]),
				.Carry_out_DO(Iteration_cell_carry_D[i])
			);
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2372:3
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2374:7
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2377:13
				if (Fsm_enable_S)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2378:16
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R1 : Iteration_cell_sum_AMASK_D[0]);
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2380:16
					Partial_remainder_DN = Partial_remainder_DP;
			2'b01:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2384:13
				if (Fsm_enable_S)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2385:16
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R2 : Iteration_cell_sum_AMASK_D[1]);
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2387:16
					Partial_remainder_DN = Partial_remainder_DP;
			2'b10:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2391:13
				if (Fsm_enable_S)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2392:16
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R3 : Iteration_cell_sum_AMASK_D[2]);
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2394:16
					Partial_remainder_DN = Partial_remainder_DP;
			2'b11:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2398:13
				if (Fsm_enable_S)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2399:16
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R4 : Iteration_cell_sum_AMASK_D[3]);
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2401:16
					Partial_remainder_DN = Partial_remainder_DP;
		endcase
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2408:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2410:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2412:14
			Partial_remainder_DP <= 1'sb0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2416:14
			Partial_remainder_DP <= Partial_remainder_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2420:4
	reg [56:0] Quotient_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2422:3
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2424:7
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2427:13
				if (Fsm_enable_S)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2428:16
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[55:0], Sqrt_quotinent_S[3]} : {Quotient_DP[55:0], Iteration_cell_carry_D[0]});
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2430:16
					Quotient_DN = Quotient_DP;
			2'b01:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2434:13
				if (Fsm_enable_S)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2435:16
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[54:0], Sqrt_quotinent_S[3:2]} : {Quotient_DP[54:0], Iteration_cell_carry_D[0], Iteration_cell_carry_D[1]});
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2437:16
					Quotient_DN = Quotient_DP;
			2'b10:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2441:13
				if (Fsm_enable_S)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2442:16
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[53:0], Sqrt_quotinent_S[3:1]} : {Quotient_DP[53:0], Iteration_cell_carry_D[0], Iteration_cell_carry_D[1], Iteration_cell_carry_D[2]});
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2444:16
					Quotient_DN = Quotient_DP;
			2'b11:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2448:13
				if (Fsm_enable_S)
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2449:16
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[defs_div_sqrt_mvp_C_MANT_FP64:0], Sqrt_quotinent_S} : {Quotient_DP[defs_div_sqrt_mvp_C_MANT_FP64:0], Iteration_cell_carry_D[0], Iteration_cell_carry_D[1], Iteration_cell_carry_D[2], Iteration_cell_carry_D[3]});
				else
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2451:16
					Quotient_DN = Quotient_DP;
		endcase
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2456:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2458:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2460:11
			Quotient_DP <= 1'sb0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2463:11
			Quotient_DP <= Quotient_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2473:4
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2814:4
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3030:4
	generate
		if (1) begin : genblk7
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3033:9
			always @(*)
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3035:13
				case (Format_sel_S)
					2'b00:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3038:19
						case (Precision_ctl_S)
							6'h00:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3041:25
								Mant_result_prenorm_DO = {Quotient_DP[26:0], {30 {1'b0}}};
							6'h17, 6'h16, 6'h15:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3045:25
								Mant_result_prenorm_DO = {Quotient_DP[defs_div_sqrt_mvp_C_MANT_FP32:0], {33 {1'b0}}};
							6'h14, 6'h13, 6'h12:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3049:25
								Mant_result_prenorm_DO = {Quotient_DP[20:0], {36 {1'b0}}};
							6'h11, 6'h10, 6'h0f:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3053:25
								Mant_result_prenorm_DO = {Quotient_DP[17:0], {39 {1'b0}}};
							6'h0e, 6'h0d, 6'h0c:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3057:25
								Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
							6'h0b, 6'h0a, 6'h09:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3061:25
								Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
							6'h08, 6'h07, 6'h06:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3065:25
								Mant_result_prenorm_DO = {Quotient_DP[8:0], {48 {1'b0}}};
							default:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3069:25
								Mant_result_prenorm_DO = {Quotient_DP[26:0], {30 {1'b0}}};
						endcase
					2'b01:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3076:19
						case (Precision_ctl_S)
							6'h00:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3079:25
								Mant_result_prenorm_DO = Quotient_DP[56:0];
							6'h34, 6'h33:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3083:25
								Mant_result_prenorm_DO = {Quotient_DP[53:1], {4 {1'b0}}};
							6'h32, 6'h31, 6'h30:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3087:25
								Mant_result_prenorm_DO = {Quotient_DP[50:0], {6 {1'b0}}};
							6'h2f, 6'h2e, 6'h2d:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3091:25
								Mant_result_prenorm_DO = {Quotient_DP[47:0], {9 {1'b0}}};
							6'h2c, 6'h2b, 6'h2a:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3095:25
								Mant_result_prenorm_DO = {Quotient_DP[44:0], {12 {1'b0}}};
							6'h29, 6'h28, 6'h27:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3099:25
								Mant_result_prenorm_DO = {Quotient_DP[41:0], {15 {1'b0}}};
							6'h26, 6'h25, 6'h24:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3103:25
								Mant_result_prenorm_DO = {Quotient_DP[38:0], {18 {1'b0}}};
							6'h23, 6'h22, 6'h21:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3107:25
								Mant_result_prenorm_DO = {Quotient_DP[35:0], {21 {1'b0}}};
							6'h20, 6'h1f, 6'h1e:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3111:25
								Mant_result_prenorm_DO = {Quotient_DP[32:0], {24 {1'b0}}};
							6'h1d, 6'h1c, 6'h1b:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3115:25
								Mant_result_prenorm_DO = {Quotient_DP[29:0], {27 {1'b0}}};
							6'h1a, 6'h19, 6'h18:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3119:25
								Mant_result_prenorm_DO = {Quotient_DP[26:0], {30 {1'b0}}};
							6'h17, 6'h16, 6'h15:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3123:25
								Mant_result_prenorm_DO = {Quotient_DP[23:0], {33 {1'b0}}};
							6'h14, 6'h13, 6'h12:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3127:25
								Mant_result_prenorm_DO = {Quotient_DP[20:0], {36 {1'b0}}};
							6'h11, 6'h10, 6'h0f:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3131:25
								Mant_result_prenorm_DO = {Quotient_DP[17:0], {39 {1'b0}}};
							6'h0e, 6'h0d, 6'h0c:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3135:25
								Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
							6'h0b, 6'h0a, 6'h09:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3139:25
								Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
							6'h08, 6'h07, 6'h06:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3143:25
								Mant_result_prenorm_DO = {Quotient_DP[8:0], {48 {1'b0}}};
							default:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3147:25
								Mant_result_prenorm_DO = Quotient_DP[56:0];
						endcase
					2'b10:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3154:19
						case (Precision_ctl_S)
							6'b000000:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3157:25
								Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
							6'h0a, 6'h09:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3161:25
								Mant_result_prenorm_DO = {Quotient_DP[11:1], {46 {1'b0}}};
							6'h08, 6'h07, 6'h06:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3165:25
								Mant_result_prenorm_DO = {Quotient_DP[8:0], {48 {1'b0}}};
							default:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3169:25
								Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
						endcase
					2'b11:
						// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3177:19
						case (Precision_ctl_S)
							6'b000000:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3180:25
								Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
							6'h07, 6'h06:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3184:25
								Mant_result_prenorm_DO = {Quotient_DP[8:1], {49 {1'b0}}};
							default:
								// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3188:25
								Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
						endcase
				endcase
		end
	endgenerate
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3199:4
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3356:4
	wire [12:0] Exp_result_prenorm_DN;
	reg [12:0] Exp_result_prenorm_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3358:4
	wire [12:0] Exp_add_a_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3359:4
	wire [12:0] Exp_add_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3360:4
	wire [12:0] Exp_add_c_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3362:3
	integer C_BIAS_AONE;
	integer C_HALF_BIAS;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3363:3
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP16 = 5'h10;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP16ALT = 8'h80;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP32 = 8'h80;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP64 = 11'h400;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP16 = 7;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP16ALT = 63;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP32 = 63;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP64 = 511;
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3365:7
		case (Format_sel_S)
			2'b00: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3368:13
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP32;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3369:13
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP32;
			end
			2'b01: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3373:13
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP64;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3374:13
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP64;
			end
			2'b10: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3378:13
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP16;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3379:13
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP16;
			end
			2'b11: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3383:13
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP16ALT;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3384:13
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP16ALT;
			end
		endcase
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3393:3
	assign Exp_add_a_D = {(Sqrt_start_dly_S ? {Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64:1]} : {Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI})};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3394:3
	localparam defs_div_sqrt_mvp_C_EXP_ZERO_FP64 = 11'h000;
	assign Exp_add_b_D = {(Sqrt_start_dly_S ? {1'b0, defs_div_sqrt_mvp_C_EXP_ZERO_FP64, Exp_num_DI[0]} : {~Exp_den_DI[defs_div_sqrt_mvp_C_EXP_FP64], ~Exp_den_DI[defs_div_sqrt_mvp_C_EXP_FP64], ~Exp_den_DI})};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3395:3
	assign Exp_add_c_D = {(Div_start_dly_S ? {C_BIAS_AONE} : {C_HALF_BIAS})};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3396:3
	assign Exp_result_prenorm_DN = (Start_dly_S ? {(Exp_add_a_D + Exp_add_b_D) + Exp_add_c_D} : Exp_result_prenorm_DP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3399:3
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3401:7
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3403:11
			Exp_result_prenorm_DP <= 1'sb0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3407:11
			Exp_result_prenorm_DP <= Exp_result_prenorm_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3411:3
	assign Exp_result_prenorm_DO = Exp_result_prenorm_DP;
endmodule
// removed package "defs_div_sqrt_mvp"
// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:44:1
// removed ["import defs_div_sqrt_mvp::*;"]
module norm_div_sqrt_mvp (
	Mant_in_DI,
	Exp_in_DI,
	Sign_in_DI,
	Div_enable_SI,
	Sqrt_enable_SI,
	Inf_a_SI,
	Inf_b_SI,
	Zero_a_SI,
	Zero_b_SI,
	NaN_a_SI,
	NaN_b_SI,
	SNaN_SI,
	RM_SI,
	Full_precision_SI,
	FP32_SI,
	FP64_SI,
	FP16_SI,
	FP16ALT_SI,
	Result_DO,
	Fflags_SO
);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:48:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	input wire [56:0] Mant_in_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:49:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	input wire signed [12:0] Exp_in_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:50:4
	input wire Sign_in_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:51:4
	input wire Div_enable_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:52:4
	input wire Sqrt_enable_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:53:4
	input wire Inf_a_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:54:4
	input wire Inf_b_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:55:4
	input wire Zero_a_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:56:4
	input wire Zero_b_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:57:4
	input wire NaN_a_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:58:4
	input wire NaN_b_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:59:4
	input wire SNaN_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:60:4
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:61:4
	input wire Full_precision_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:62:4
	input wire FP32_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:63:4
	input wire FP64_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:64:4
	input wire FP16_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:65:4
	input wire FP16ALT_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:67:4
	output reg [63:0] Result_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:68:4
	output wire [4:0] Fflags_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:72:4
	reg Sign_res_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:74:4
	reg NV_OP_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:75:4
	reg Exp_OF_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:76:4
	reg Exp_UF_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:77:4
	reg Div_Zero_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:78:4
	wire In_Exact_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:83:4
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_res_norm_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:84:4
	reg [10:0] Exp_res_norm_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:90:3
	wire [12:0] Exp_Max_RS_FP64_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:91:3
	localparam defs_div_sqrt_mvp_C_EXP_FP32 = 8;
	wire [9:0] Exp_Max_RS_FP32_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:92:3
	localparam defs_div_sqrt_mvp_C_EXP_FP16 = 5;
	wire [6:0] Exp_Max_RS_FP16_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:93:3
	localparam defs_div_sqrt_mvp_C_EXP_FP16ALT = 8;
	wire [9:0] Exp_Max_RS_FP16ALT_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:95:3
	assign Exp_Max_RS_FP64_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64:0] + defs_div_sqrt_mvp_C_MANT_FP64) + 1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:96:3
	localparam defs_div_sqrt_mvp_C_MANT_FP32 = 23;
	assign Exp_Max_RS_FP32_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP32:0] + defs_div_sqrt_mvp_C_MANT_FP32) + 1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:97:3
	localparam defs_div_sqrt_mvp_C_MANT_FP16 = 10;
	assign Exp_Max_RS_FP16_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16:0] + defs_div_sqrt_mvp_C_MANT_FP16) + 1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:98:3
	localparam defs_div_sqrt_mvp_C_MANT_FP16ALT = 7;
	assign Exp_Max_RS_FP16ALT_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16ALT:0] + defs_div_sqrt_mvp_C_MANT_FP16ALT) + 1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:99:3
	wire [12:0] Num_RS_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:100:3
	assign Num_RS_D = ~Exp_in_DI + 2;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:101:3
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_RS_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:102:3
	wire [56:0] Mant_forsticky_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:103:3
	assign {Mant_RS_D, Mant_forsticky_D} = {Mant_in_DI, {53 {1'b0}}} >> Num_RS_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:105:3
	wire [12:0] Exp_subOne_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:106:3
	assign Exp_subOne_D = Exp_in_DI - 1;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:109:4
	reg [1:0] Mant_lower_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:110:4
	reg Mant_sticky_bit_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:111:4
	reg [56:0] Mant_forround_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:113:4
	localparam defs_div_sqrt_mvp_C_EXP_ONE_FP64 = 13'h0001;
	localparam defs_div_sqrt_mvp_C_MANT_NAN_FP64 = 52'h8000000000000;
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:116:8
		if (NaN_a_SI) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:118:12
			Div_Zero_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:119:12
			Exp_OF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:120:12
			Exp_UF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:121:12
			Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:122:12
			Exp_res_norm_D = 1'sb1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:123:12
			Mant_forround_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:124:12
			Sign_res_D = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:125:12
			NV_OP_S = SNaN_SI;
		end
		else if (NaN_b_SI) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:130:11
			Div_Zero_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:131:11
			Exp_OF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:132:11
			Exp_UF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:133:11
			Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:134:11
			Exp_res_norm_D = 1'sb1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:135:11
			Mant_forround_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:136:11
			Sign_res_D = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:137:11
			NV_OP_S = SNaN_SI;
		end
		else if (Inf_a_SI) begin
			begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:142:11
				if (Div_enable_SI && Inf_b_SI) begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:144:15
					Div_Zero_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:145:15
					Exp_OF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:146:15
					Exp_UF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:147:15
					Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:148:15
					Exp_res_norm_D = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:149:15
					Mant_forround_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:150:15
					Sign_res_D = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:151:15
					NV_OP_S = 1'b1;
				end
				else if (Sqrt_enable_SI && Sign_in_DI) begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:154:13
					Div_Zero_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:155:13
					Exp_OF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:156:13
					Exp_UF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:157:13
					Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:158:13
					Exp_res_norm_D = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:159:13
					Mant_forround_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:160:13
					Sign_res_D = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:161:13
					NV_OP_S = 1'b1;
				end
				else begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:163:13
					Div_Zero_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:164:13
					Exp_OF_S = 1'b1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:165:13
					Exp_UF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:166:13
					Mant_res_norm_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:167:13
					Exp_res_norm_D = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:168:13
					Mant_forround_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:169:13
					Sign_res_D = Sign_in_DI;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:170:13
					NV_OP_S = 1'b0;
				end
			end
		end
		else if (Div_enable_SI && Inf_b_SI) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:176:11
			Div_Zero_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:177:11
			Exp_OF_S = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:178:11
			Exp_UF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:179:11
			Mant_res_norm_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:180:11
			Exp_res_norm_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:181:11
			Mant_forround_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:182:11
			Sign_res_D = Sign_in_DI;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:183:11
			NV_OP_S = 1'b0;
		end
		else if (Zero_a_SI) begin
			begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:188:10
				if (Div_enable_SI && Zero_b_SI) begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:190:15
					Div_Zero_S = 1'b1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:191:15
					Exp_OF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:192:15
					Exp_UF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:193:15
					Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:194:15
					Exp_res_norm_D = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:195:15
					Mant_forround_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:196:15
					Sign_res_D = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:197:15
					NV_OP_S = 1'b1;
				end
				else begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:201:14
					Div_Zero_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:202:14
					Exp_OF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:203:14
					Exp_UF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:204:14
					Mant_res_norm_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:205:14
					Exp_res_norm_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:206:14
					Mant_forround_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:207:14
					Sign_res_D = Sign_in_DI;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:208:14
					NV_OP_S = 1'b0;
				end
			end
		end
		else if (Div_enable_SI && Zero_b_SI) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:214:10
			Div_Zero_S = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:215:10
			Exp_OF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:216:10
			Exp_UF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:217:10
			Mant_res_norm_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:218:10
			Exp_res_norm_D = 1'sb1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:219:10
			Mant_forround_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:220:10
			Sign_res_D = Sign_in_DI;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:221:10
			NV_OP_S = 1'b0;
		end
		else if (Sign_in_DI && Sqrt_enable_SI) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:226:11
			Div_Zero_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:227:11
			Exp_OF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:228:11
			Exp_UF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:229:11
			Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:230:11
			Exp_res_norm_D = 1'sb1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:231:11
			Mant_forround_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:232:11
			Sign_res_D = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:233:11
			NV_OP_S = 1'b1;
		end
		else if (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64:0] == {12 {1'sb0}}) begin
			begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:238:10
				if (Mant_in_DI != {57 {1'sb0}}) begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:240:14
					Div_Zero_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:241:14
					Exp_OF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:242:14
					Exp_UF_S = 1'b1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:243:14
					Mant_res_norm_D = {1'b0, Mant_in_DI[56:5]};
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:244:14
					Exp_res_norm_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:245:14
					Mant_forround_D = {Mant_in_DI[4:0], {defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}};
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:246:14
					Sign_res_D = Sign_in_DI;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:247:14
					NV_OP_S = 1'b0;
				end
				else begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:251:14
					Div_Zero_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:252:14
					Exp_OF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:253:14
					Exp_UF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:254:14
					Mant_res_norm_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:255:14
					Exp_res_norm_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:256:14
					Mant_forround_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:257:14
					Sign_res_D = Sign_in_DI;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:258:14
					NV_OP_S = 1'b0;
				end
			end
		end
		else if ((Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64:0] == defs_div_sqrt_mvp_C_EXP_ONE_FP64) && ~Mant_in_DI[56]) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:264:11
			Div_Zero_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:265:11
			Exp_OF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:266:11
			Exp_UF_S = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:267:11
			Mant_res_norm_D = Mant_in_DI[56:4];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:268:11
			Exp_res_norm_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:269:11
			Mant_forround_D = {Mant_in_DI[3:0], {53 {1'b0}}};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:270:11
			Sign_res_D = Sign_in_DI;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:271:11
			NV_OP_S = 1'b0;
		end
		else if (Exp_in_DI[12]) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:276:11
			Div_Zero_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:277:11
			Exp_OF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:278:11
			Exp_UF_S = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:279:11
			Mant_res_norm_D = {Mant_RS_D[defs_div_sqrt_mvp_C_MANT_FP64:0]};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:280:11
			Exp_res_norm_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:281:11
			Mant_forround_D = {Mant_forsticky_D[56:0]};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:282:11
			Sign_res_D = Sign_in_DI;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:283:11
			NV_OP_S = 1'b0;
		end
		else if ((((Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP32] && FP32_SI) | (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64] && FP64_SI)) | (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16] && FP16_SI)) | (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16ALT] && FP16ALT_SI)) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:288:11
			Div_Zero_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:289:11
			Exp_OF_S = 1'b1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:290:11
			Exp_UF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:291:11
			Mant_res_norm_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:292:11
			Exp_res_norm_D = 1'sb1;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:293:11
			Mant_forround_D = 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:294:11
			Sign_res_D = Sign_in_DI;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:295:11
			NV_OP_S = 1'b0;
		end
		else if (((((Exp_in_DI[7:0] == {8 {1'sb1}}) && FP32_SI) | ((Exp_in_DI[10:0] == {11 {1'sb1}}) && FP64_SI)) | ((Exp_in_DI[4:0] == {5 {1'sb1}}) && FP16_SI)) | ((Exp_in_DI[7:0] == {8 {1'sb1}}) && FP16ALT_SI)) begin
			begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:300:11
				if (~Mant_in_DI[56]) begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:302:15
					Div_Zero_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:303:15
					Exp_OF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:304:15
					Exp_UF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:305:15
					Mant_res_norm_D = Mant_in_DI[55:3];
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:306:15
					Exp_res_norm_D = Exp_subOne_D;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:307:15
					Mant_forround_D = {Mant_in_DI[2:0], {54 {1'b0}}};
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:308:15
					Sign_res_D = Sign_in_DI;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:309:15
					NV_OP_S = 1'b0;
				end
				else if (Mant_in_DI != {57 {1'sb0}}) begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:313:15
					Div_Zero_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:314:15
					Exp_OF_S = 1'b1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:315:15
					Exp_UF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:316:15
					Mant_res_norm_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:317:15
					Exp_res_norm_D = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:318:15
					Mant_forround_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:319:15
					Sign_res_D = Sign_in_DI;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:320:15
					NV_OP_S = 1'b0;
				end
				else begin
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:324:15
					Div_Zero_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:325:15
					Exp_OF_S = 1'b1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:326:15
					Exp_UF_S = 1'b0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:327:15
					Mant_res_norm_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:328:15
					Exp_res_norm_D = 1'sb1;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:329:15
					Mant_forround_D = 1'sb0;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:330:15
					Sign_res_D = Sign_in_DI;
					// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:331:15
					NV_OP_S = 1'b0;
				end
			end
		end
		else if (Mant_in_DI[56]) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:337:12
			Div_Zero_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:338:12
			Exp_OF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:339:12
			Exp_UF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:340:12
			Mant_res_norm_D = Mant_in_DI[56:4];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:341:12
			Exp_res_norm_D = Exp_in_DI[10:0];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:342:12
			Mant_forround_D = {Mant_in_DI[3:0], {53 {1'b0}}};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:343:12
			Sign_res_D = Sign_in_DI;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:344:12
			NV_OP_S = 1'b0;
		end
		else begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:349:12
			Div_Zero_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:350:12
			Exp_OF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:351:12
			Exp_UF_S = 1'b0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:352:12
			Mant_res_norm_D = Mant_in_DI[55:3];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:353:12
			Exp_res_norm_D = Exp_subOne_D;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:354:12
			Mant_forround_D = {Mant_in_DI[2:0], {54 {1'b0}}};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:355:12
			Sign_res_D = Sign_in_DI;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:356:12
			NV_OP_S = 1'b0;
		end
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:365:4
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_upper_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:366:4
	wire [53:0] Mant_upperRounded_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:367:4
	reg Mant_roundUp_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:368:4
	wire Mant_rounded_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:370:3
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:372:7
		if (FP32_SI) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:374:11
			Mant_upper_D = {Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:29], {29 {1'b0}}};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:375:11
			Mant_lower_D = Mant_res_norm_D[28:27];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:376:11
			Mant_sticky_bit_D = |Mant_res_norm_D[26:0];
		end
		else if (FP64_SI) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:380:11
			Mant_upper_D = Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:0];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:381:11
			Mant_lower_D = Mant_forround_D[56:55];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:382:11
			Mant_sticky_bit_D = |Mant_forround_D[55:0];
		end
		else if (FP16_SI) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:386:11
			Mant_upper_D = {Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:42], {42 {1'b0}}};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:387:11
			Mant_lower_D = Mant_res_norm_D[41:40];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:388:11
			Mant_sticky_bit_D = |Mant_res_norm_D[39:30];
		end
		else begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:392:11
			Mant_upper_D = {Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:45], {45 {1'b0}}};
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:393:11
			Mant_lower_D = Mant_res_norm_D[44:43];
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:394:11
			Mant_sticky_bit_D = |Mant_res_norm_D[42:30];
		end
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:398:4
	assign Mant_rounded_S = |Mant_lower_D | Mant_sticky_bit_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:403:4
	localparam defs_div_sqrt_mvp_C_RM_MINUSINF = 3'h3;
	localparam defs_div_sqrt_mvp_C_RM_NEAREST = 3'h0;
	localparam defs_div_sqrt_mvp_C_RM_PLUSINF = 3'h2;
	localparam defs_div_sqrt_mvp_C_RM_TRUNC = 3'h1;
	always @(*) begin
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:405:9
		Mant_roundUp_S = 1'b0;
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:406:9
		case (RM_SI)
			defs_div_sqrt_mvp_C_RM_NEAREST:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:408:13
				Mant_roundUp_S = Mant_lower_D[1] && ((Mant_lower_D[0] | Mant_sticky_bit_D) | ((((FP32_SI && Mant_upper_D[29]) | (FP64_SI && Mant_upper_D[0])) | (FP16_SI && Mant_upper_D[42])) | (FP16ALT_SI && Mant_upper_D[45])));
			defs_div_sqrt_mvp_C_RM_TRUNC:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:410:13
				Mant_roundUp_S = 0;
			defs_div_sqrt_mvp_C_RM_PLUSINF:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:412:13
				Mant_roundUp_S = Mant_rounded_S & ~Sign_in_DI;
			defs_div_sqrt_mvp_C_RM_MINUSINF:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:414:13
				Mant_roundUp_S = Mant_rounded_S & Sign_in_DI;
			default:
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:416:13
				Mant_roundUp_S = 0;
		endcase
	end
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:420:3
	wire Mant_renorm_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:421:3
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_roundUp_Vector_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:423:3
	assign Mant_roundUp_Vector_S = {7'h00, FP16ALT_SI && Mant_roundUp_S, 2'h0, FP16_SI && Mant_roundUp_S, 12'h000, FP32_SI && Mant_roundUp_S, 28'h0000000, FP64_SI && Mant_roundUp_S};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:426:3
	assign Mant_upperRounded_D = Mant_upper_D + Mant_roundUp_Vector_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:427:3
	assign Mant_renorm_S = Mant_upperRounded_D[53];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:432:3
	wire [51:0] Mant_res_round_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:433:3
	wire [10:0] Exp_res_round_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:436:3
	assign Mant_res_round_D = (Mant_renorm_S ? Mant_upperRounded_D[defs_div_sqrt_mvp_C_MANT_FP64:1] : Mant_upperRounded_D[51:0]);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:437:3
	assign Exp_res_round_D = Exp_res_norm_D + Mant_renorm_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:442:3
	wire [51:0] Mant_before_format_ctl_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:443:3
	wire [10:0] Exp_before_format_ctl_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:444:3
	assign Mant_before_format_ctl_D = (Full_precision_SI ? Mant_res_round_D : Mant_res_norm_D);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:445:3
	assign Exp_before_format_ctl_D = (Full_precision_SI ? Exp_res_round_D : Exp_res_norm_D);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:447:3
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:449:7
		if (FP32_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:451:13
			Result_DO = {32'hffffffff, Sign_res_D, Exp_before_format_ctl_D[7:0], Mant_before_format_ctl_D[51:29]};
		else if (FP64_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:455:13
			Result_DO = {Sign_res_D, Exp_before_format_ctl_D[10:0], Mant_before_format_ctl_D[51:0]};
		else if (FP16_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:459:13
			Result_DO = {48'hffffffffffff, Sign_res_D, Exp_before_format_ctl_D[4:0], Mant_before_format_ctl_D[51:42]};
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:463:13
			Result_DO = {48'hffffffffffff, Sign_res_D, Exp_before_format_ctl_D[7:0], Mant_before_format_ctl_D[51:45]};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:467:1
	assign In_Exact_S = ~Full_precision_SI | Mant_rounded_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:468:1
	assign Fflags_SO = {NV_OP_S, Div_Zero_S, Exp_OF_S, Exp_UF_S, In_Exact_S};
endmodule
// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:34:1
// removed ["import defs_div_sqrt_mvp::*;"]
module nrbd_nrsc_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Start_SI,
	Kill_SI,
	Special_case_SBI,
	Special_case_dly_SBI,
	Precision_ctl_SI,
	Format_sel_SI,
	Mant_a_DI,
	Mant_b_DI,
	Exp_a_DI,
	Exp_b_DI,
	Div_enable_SO,
	Sqrt_enable_SO,
	Full_precision_SO,
	FP32_SO,
	FP64_SO,
	FP16_SO,
	FP16ALT_SO,
	Ready_SO,
	Done_SO,
	Mant_z_DO,
	Exp_z_DO
);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:39:4
	input wire Clk_CI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:40:4
	input wire Rst_RBI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:41:4
	input wire Div_start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:42:4
	input wire Sqrt_start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:43:4
	input wire Start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:44:4
	input wire Kill_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:45:4
	input wire Special_case_SBI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:46:4
	input wire Special_case_dly_SBI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:47:4
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:48:4
	input wire [1:0] Format_sel_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:49:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:50:4
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:51:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:52:4
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:54:4
	output wire Div_enable_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:55:4
	output wire Sqrt_enable_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:57:4
	output wire Full_precision_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:58:4
	output wire FP32_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:59:4
	output wire FP64_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:60:4
	output wire FP16_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:61:4
	output wire FP16ALT_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:62:4
	output wire Ready_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:63:4
	output wire Done_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:64:4
	output wire [56:0] Mant_z_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:65:4
	output wire [12:0] Exp_z_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:69:5
	wire Div_start_dly_S;
	wire Sqrt_start_dly_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:72:1
	control_mvp control_U0(
		.Clk_CI(Clk_CI),
		.Rst_RBI(Rst_RBI),
		.Div_start_SI(Div_start_SI),
		.Sqrt_start_SI(Sqrt_start_SI),
		.Start_SI(Start_SI),
		.Kill_SI(Kill_SI),
		.Special_case_SBI(Special_case_SBI),
		.Special_case_dly_SBI(Special_case_dly_SBI),
		.Precision_ctl_SI(Precision_ctl_SI),
		.Format_sel_SI(Format_sel_SI),
		.Numerator_DI(Mant_a_DI),
		.Exp_num_DI(Exp_a_DI),
		.Denominator_DI(Mant_b_DI),
		.Exp_den_DI(Exp_b_DI),
		.Div_start_dly_SO(Div_start_dly_S),
		.Sqrt_start_dly_SO(Sqrt_start_dly_S),
		.Div_enable_SO(Div_enable_SO),
		.Sqrt_enable_SO(Sqrt_enable_SO),
		.Full_precision_SO(Full_precision_SO),
		.FP32_SO(FP32_SO),
		.FP64_SO(FP64_SO),
		.FP16_SO(FP16_SO),
		.FP16ALT_SO(FP16ALT_SO),
		.Ready_SO(Ready_SO),
		.Done_SO(Done_SO),
		.Mant_result_prenorm_DO(Mant_z_DO),
		.Exp_result_prenorm_DO(Exp_z_DO)
	);
endmodule
module iteration_div_sqrt_mvp (
	A_DI,
	B_DI,
	Div_enable_SI,
	Div_start_dly_SI,
	Sqrt_enable_SI,
	D_DI,
	D_DO,
	Sum_DO,
	Carry_out_DO
);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:34:16
	parameter WIDTH = 25;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:38:4
	input wire [WIDTH - 1:0] A_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:39:4
	input wire [WIDTH - 1:0] B_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:40:4
	input wire Div_enable_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:41:4
	input wire Div_start_dly_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:42:4
	input wire Sqrt_enable_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:43:4
	input wire [1:0] D_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:45:4
	output wire [1:0] D_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:46:4
	output wire [WIDTH - 1:0] Sum_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:47:4
	output wire Carry_out_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:50:4
	wire D_carry_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:51:4
	wire Sqrt_cin_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:52:4
	wire Cin_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:54:4
	assign D_DO[0] = ~D_DI[0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:55:4
	assign D_DO[1] = ~(D_DI[1] ^ D_DI[0]);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:56:4
	assign D_carry_D = D_DI[1] | D_DI[0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:57:4
	assign Sqrt_cin_D = Sqrt_enable_SI && D_carry_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:58:4
	assign Cin_D = (Div_enable_SI ? 1'b0 : Sqrt_cin_D);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:59:4
	assign {Carry_out_DO, Sum_DO} = (A_DI + B_DI) + Cin_D;
endmodule
// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:35:1
// removed ["import defs_div_sqrt_mvp::*;"]
module div_sqrt_top_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Operand_a_DI,
	Operand_b_DI,
	RM_SI,
	Precision_ctl_SI,
	Format_sel_SI,
	Kill_SI,
	Result_DO,
	Fflags_SO,
	Ready_SO,
	Done_SO
);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:40:4
	input wire Clk_CI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:41:4
	input wire Rst_RBI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:42:4
	input wire Div_start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:43:4
	input wire Sqrt_start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:46:4
	localparam defs_div_sqrt_mvp_C_OP_FP64 = 64;
	input wire [63:0] Operand_a_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:47:4
	input wire [63:0] Operand_b_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:50:4
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:51:4
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:52:4
	localparam defs_div_sqrt_mvp_C_FS = 2;
	input wire [1:0] Format_sel_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:53:4
	input wire Kill_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:56:4
	output wire [63:0] Result_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:59:4
	output wire [4:0] Fflags_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:60:4
	output wire Ready_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:61:4
	output wire Done_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:69:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:70:4
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:71:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:72:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:74:4
	wire [12:0] Exp_z_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:75:4
	wire [56:0] Mant_z_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:76:4
	wire Sign_z_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:77:4
	wire Start_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:78:4
	wire [2:0] RM_dly_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:79:4
	wire Div_enable_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:80:4
	wire Sqrt_enable_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:81:4
	wire Inf_a_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:82:4
	wire Inf_b_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:83:4
	wire Zero_a_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:84:4
	wire Zero_b_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:85:4
	wire NaN_a_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:86:4
	wire NaN_b_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:87:4
	wire SNaN_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:88:4
	wire Special_case_SB;
	wire Special_case_dly_SB;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:90:4
	wire Full_precision_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:91:4
	wire FP32_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:92:4
	wire FP64_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:93:4
	wire FP16_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:94:4
	wire FP16ALT_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:97:2
	preprocess_mvp preprocess_U0(
		.Clk_CI(Clk_CI),
		.Rst_RBI(Rst_RBI),
		.Div_start_SI(Div_start_SI),
		.Sqrt_start_SI(Sqrt_start_SI),
		.Ready_SI(Ready_SO),
		.Operand_a_DI(Operand_a_DI),
		.Operand_b_DI(Operand_b_DI),
		.RM_SI(RM_SI),
		.Format_sel_SI(Format_sel_SI),
		.Start_SO(Start_S),
		.Exp_a_DO_norm(Exp_a_D),
		.Exp_b_DO_norm(Exp_b_D),
		.Mant_a_DO_norm(Mant_a_D),
		.Mant_b_DO_norm(Mant_b_D),
		.RM_dly_SO(RM_dly_S),
		.Sign_z_DO(Sign_z_D),
		.Inf_a_SO(Inf_a_S),
		.Inf_b_SO(Inf_b_S),
		.Zero_a_SO(Zero_a_S),
		.Zero_b_SO(Zero_b_S),
		.NaN_a_SO(NaN_a_S),
		.NaN_b_SO(NaN_b_S),
		.SNaN_SO(SNaN_S),
		.Special_case_SBO(Special_case_SB),
		.Special_case_dly_SBO(Special_case_dly_SB)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:126:2
	nrbd_nrsc_mvp nrbd_nrsc_U0(
		.Clk_CI(Clk_CI),
		.Rst_RBI(Rst_RBI),
		.Div_start_SI(Div_start_SI),
		.Sqrt_start_SI(Sqrt_start_SI),
		.Start_SI(Start_S),
		.Kill_SI(Kill_SI),
		.Special_case_SBI(Special_case_SB),
		.Special_case_dly_SBI(Special_case_dly_SB),
		.Div_enable_SO(Div_enable_S),
		.Sqrt_enable_SO(Sqrt_enable_S),
		.Precision_ctl_SI(Precision_ctl_SI),
		.Format_sel_SI(Format_sel_SI),
		.Exp_a_DI(Exp_a_D),
		.Exp_b_DI(Exp_b_D),
		.Mant_a_DI(Mant_a_D),
		.Mant_b_DI(Mant_b_D),
		.Full_precision_SO(Full_precision_S),
		.FP32_SO(FP32_S),
		.FP64_SO(FP64_S),
		.FP16_SO(FP16_S),
		.FP16ALT_SO(FP16ALT_S),
		.Ready_SO(Ready_SO),
		.Done_SO(Done_SO),
		.Exp_z_DO(Exp_z_D),
		.Mant_z_DO(Mant_z_D)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:156:2
	norm_div_sqrt_mvp fpu_norm_U0(
		.Mant_in_DI(Mant_z_D),
		.Exp_in_DI(Exp_z_D),
		.Sign_in_DI(Sign_z_D),
		.Div_enable_SI(Div_enable_S),
		.Sqrt_enable_SI(Sqrt_enable_S),
		.Inf_a_SI(Inf_a_S),
		.Inf_b_SI(Inf_b_S),
		.Zero_a_SI(Zero_a_S),
		.Zero_b_SI(Zero_b_S),
		.NaN_a_SI(NaN_a_S),
		.NaN_b_SI(NaN_b_S),
		.SNaN_SI(SNaN_S),
		.RM_SI(RM_dly_S),
		.Full_precision_SI(Full_precision_S),
		.FP32_SI(FP32_S),
		.FP64_SI(FP64_S),
		.FP16_SI(FP16_S),
		.FP16ALT_SI(FP16ALT_S),
		.Result_DO(Result_DO),
		.Fflags_SO(Fflags_SO)
	);
endmodule
// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:39:1
// removed ["import defs_div_sqrt_mvp::*;"]
// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:35:1
// removed ["import defs_div_sqrt_mvp::*;"]
module preprocess_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Ready_SI,
	Operand_a_DI,
	Operand_b_DI,
	RM_SI,
	Format_sel_SI,
	Start_SO,
	Exp_a_DO_norm,
	Exp_b_DO_norm,
	Mant_a_DO_norm,
	Mant_b_DO_norm,
	RM_dly_SO,
	Sign_z_DO,
	Inf_a_SO,
	Inf_b_SO,
	Zero_a_SO,
	Zero_b_SO,
	NaN_a_SO,
	NaN_b_SO,
	SNaN_SO,
	Special_case_SBO,
	Special_case_dly_SBO
);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:39:4
	input wire Clk_CI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:40:4
	input wire Rst_RBI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:41:4
	input wire Div_start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:42:4
	input wire Sqrt_start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:43:4
	input wire Ready_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:45:4
	localparam defs_div_sqrt_mvp_C_OP_FP64 = 64;
	input wire [63:0] Operand_a_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:46:4
	input wire [63:0] Operand_b_DI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:47:4
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:48:4
	localparam defs_div_sqrt_mvp_C_FS = 2;
	input wire [1:0] Format_sel_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:51:4
	output wire Start_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:52:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	output wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_DO_norm;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:53:4
	output wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_DO_norm;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:54:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	output wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_DO_norm;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:55:4
	output wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_DO_norm;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:57:4
	output wire [2:0] RM_dly_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:59:4
	output wire Sign_z_DO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:60:4
	output wire Inf_a_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:61:4
	output wire Inf_b_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:62:4
	output wire Zero_a_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:63:4
	output wire Zero_b_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:64:4
	output wire NaN_a_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:65:4
	output wire NaN_b_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:66:4
	output wire SNaN_SO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:67:4
	output wire Special_case_SBO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:68:4
	output reg Special_case_dly_SBO;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:72:4
	wire Hb_a_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:73:4
	wire Hb_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:75:4
	reg [10:0] Exp_a_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:76:4
	reg [10:0] Exp_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:77:4
	reg [51:0] Mant_a_NonH_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:78:4
	reg [51:0] Mant_b_NonH_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:79:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:80:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:85:4
	reg Sign_a_D;
	reg Sign_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:86:4
	wire Start_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:88:6
	localparam defs_div_sqrt_mvp_C_MANT_FP16 = 10;
	localparam defs_div_sqrt_mvp_C_MANT_FP16ALT = 7;
	localparam defs_div_sqrt_mvp_C_MANT_FP32 = 23;
	localparam defs_div_sqrt_mvp_C_OP_FP16 = 16;
	localparam defs_div_sqrt_mvp_C_OP_FP16ALT = 16;
	localparam defs_div_sqrt_mvp_C_OP_FP32 = 32;
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:90:10
		case (Format_sel_SI)
			2'b00: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:93:16
				Sign_a_D = Operand_a_DI[31];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:94:16
				Sign_b_D = Operand_b_DI[31];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:95:16
				Exp_a_D = {3'h0, Operand_a_DI[30:defs_div_sqrt_mvp_C_MANT_FP32]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:96:16
				Exp_b_D = {3'h0, Operand_b_DI[30:defs_div_sqrt_mvp_C_MANT_FP32]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:97:16
				Mant_a_NonH_D = {Operand_a_DI[22:0], 29'h00000000};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:98:16
				Mant_b_NonH_D = {Operand_b_DI[22:0], 29'h00000000};
			end
			2'b01: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:102:16
				Sign_a_D = Operand_a_DI[63];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:103:16
				Sign_b_D = Operand_b_DI[63];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:104:16
				Exp_a_D = Operand_a_DI[62:defs_div_sqrt_mvp_C_MANT_FP64];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:105:16
				Exp_b_D = Operand_b_DI[62:defs_div_sqrt_mvp_C_MANT_FP64];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:106:16
				Mant_a_NonH_D = Operand_a_DI[51:0];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:107:16
				Mant_b_NonH_D = Operand_b_DI[51:0];
			end
			2'b10: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:111:16
				Sign_a_D = Operand_a_DI[15];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:112:16
				Sign_b_D = Operand_b_DI[15];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:113:16
				Exp_a_D = {6'h00, Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:114:16
				Exp_b_D = {6'h00, Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:115:16
				Mant_a_NonH_D = {Operand_a_DI[9:0], 42'h00000000000};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:116:16
				Mant_b_NonH_D = {Operand_b_DI[9:0], 42'h00000000000};
			end
			2'b11: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:120:16
				Sign_a_D = Operand_a_DI[15];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:121:16
				Sign_b_D = Operand_b_DI[15];
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:122:16
				Exp_a_D = {3'h0, Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:123:16
				Exp_b_D = {3'h0, Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT]};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:124:16
				Mant_a_NonH_D = {Operand_a_DI[6:0], 45'h000000000000};
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:125:16
				Mant_b_NonH_D = {Operand_b_DI[6:0], 45'h000000000000};
			end
		endcase
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:131:4
	assign Mant_a_D = {Hb_a_D, Mant_a_NonH_D};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:132:4
	assign Mant_b_D = {Hb_b_D, Mant_b_NonH_D};
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:134:4
	assign Hb_a_D = |Exp_a_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:135:4
	assign Hb_b_D = |Exp_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:137:4
	assign Start_S = Div_start_SI | Sqrt_start_SI;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:145:4
	reg Mant_a_prenorm_zero_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:146:4
	reg Mant_b_prenorm_zero_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:148:4
	wire Exp_a_prenorm_zero_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:149:4
	wire Exp_b_prenorm_zero_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:150:4
	assign Exp_a_prenorm_zero_S = ~Hb_a_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:151:4
	assign Exp_b_prenorm_zero_S = ~Hb_b_D;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:153:4
	reg Exp_a_prenorm_Inf_NaN_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:154:4
	reg Exp_b_prenorm_Inf_NaN_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:156:4
	wire Mant_a_prenorm_QNaN_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:157:4
	wire Mant_a_prenorm_SNaN_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:158:4
	wire Mant_b_prenorm_QNaN_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:159:4
	wire Mant_b_prenorm_SNaN_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:161:4
	assign Mant_a_prenorm_QNaN_S = Mant_a_NonH_D[51] && ~(|Mant_a_NonH_D[50:0]);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:162:4
	assign Mant_a_prenorm_SNaN_S = ~Mant_a_NonH_D[51] && |Mant_a_NonH_D[50:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:163:4
	assign Mant_b_prenorm_QNaN_S = Mant_b_NonH_D[51] && ~(|Mant_b_NonH_D[50:0]);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:164:4
	assign Mant_b_prenorm_SNaN_S = ~Mant_b_NonH_D[51] && |Mant_b_NonH_D[50:0];
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:166:6
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP16 = 5'h1f;
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP16ALT = 8'hff;
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP32 = 8'hff;
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP64 = 11'h7ff;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP16 = 10'h000;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP16ALT = 7'h00;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP32 = 23'h000000;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP64 = 52'h0000000000000;
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:168:10
		case (Format_sel_SI)
			2'b00: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:171:16
				Mant_a_prenorm_zero_S = Operand_a_DI[22:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP32;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:172:16
				Mant_b_prenorm_zero_S = Operand_b_DI[22:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP32;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:173:16
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[30:defs_div_sqrt_mvp_C_MANT_FP32] == defs_div_sqrt_mvp_C_EXP_INF_FP32;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:174:16
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[30:defs_div_sqrt_mvp_C_MANT_FP32] == defs_div_sqrt_mvp_C_EXP_INF_FP32;
			end
			2'b01: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:178:16
				Mant_a_prenorm_zero_S = Operand_a_DI[51:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP64;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:179:16
				Mant_b_prenorm_zero_S = Operand_b_DI[51:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP64;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:180:16
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[62:defs_div_sqrt_mvp_C_MANT_FP64] == defs_div_sqrt_mvp_C_EXP_INF_FP64;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:181:16
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[62:defs_div_sqrt_mvp_C_MANT_FP64] == defs_div_sqrt_mvp_C_EXP_INF_FP64;
			end
			2'b10: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:185:16
				Mant_a_prenorm_zero_S = Operand_a_DI[9:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:186:16
				Mant_b_prenorm_zero_S = Operand_b_DI[9:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:187:16
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16] == defs_div_sqrt_mvp_C_EXP_INF_FP16;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:188:16
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16] == defs_div_sqrt_mvp_C_EXP_INF_FP16;
			end
			2'b11: begin
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:192:16
				Mant_a_prenorm_zero_S = Operand_a_DI[6:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16ALT;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:193:16
				Mant_b_prenorm_zero_S = Operand_b_DI[6:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16ALT;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:194:16
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT] == defs_div_sqrt_mvp_C_EXP_INF_FP16ALT;
				// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:195:16
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT] == defs_div_sqrt_mvp_C_EXP_INF_FP16ALT;
			end
		endcase
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:203:4
	wire Zero_a_SN;
	reg Zero_a_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:204:4
	wire Zero_b_SN;
	reg Zero_b_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:205:4
	wire Inf_a_SN;
	reg Inf_a_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:206:4
	wire Inf_b_SN;
	reg Inf_b_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:207:4
	wire NaN_a_SN;
	reg NaN_a_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:208:4
	wire NaN_b_SN;
	reg NaN_b_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:209:4
	wire SNaN_SN;
	reg SNaN_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:211:4
	assign Zero_a_SN = (Start_S && Ready_SI ? Exp_a_prenorm_zero_S && Mant_a_prenorm_zero_S : Zero_a_SP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:212:4
	assign Zero_b_SN = (Start_S && Ready_SI ? Exp_b_prenorm_zero_S && Mant_b_prenorm_zero_S : Zero_b_SP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:213:4
	assign Inf_a_SN = (Start_S && Ready_SI ? Exp_a_prenorm_Inf_NaN_S && Mant_a_prenorm_zero_S : Inf_a_SP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:214:4
	assign Inf_b_SN = (Start_S && Ready_SI ? Exp_b_prenorm_Inf_NaN_S && Mant_b_prenorm_zero_S : Inf_b_SP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:215:4
	assign NaN_a_SN = (Start_S && Ready_SI ? Exp_a_prenorm_Inf_NaN_S && ~Mant_a_prenorm_zero_S : NaN_a_SP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:216:4
	assign NaN_b_SN = (Start_S && Ready_SI ? Exp_b_prenorm_Inf_NaN_S && ~Mant_b_prenorm_zero_S : NaN_b_SP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:217:4
	assign SNaN_SN = (Start_S && Ready_SI ? (Mant_a_prenorm_SNaN_S && NaN_a_SN) | (Mant_b_prenorm_SNaN_S && NaN_b_SN) : SNaN_SP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:219:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:221:9
		if (~Rst_RBI) begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:223:13
			Zero_a_SP <= 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:224:13
			Zero_b_SP <= 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:225:13
			Inf_a_SP <= 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:226:13
			Inf_b_SP <= 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:227:13
			NaN_a_SP <= 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:228:13
			NaN_b_SP <= 1'sb0;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:229:13
			SNaN_SP <= 1'sb0;
		end
		else begin
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:233:12
			Inf_a_SP <= Inf_a_SN;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:234:12
			Inf_b_SP <= Inf_b_SN;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:235:12
			Zero_a_SP <= Zero_a_SN;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:236:12
			Zero_b_SP <= Zero_b_SN;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:237:12
			NaN_a_SP <= NaN_a_SN;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:238:12
			NaN_b_SP <= NaN_b_SN;
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:239:12
			SNaN_SP <= SNaN_SN;
		end
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:247:4
	assign Special_case_SBO = ~{(Div_start_SI ? ((((Zero_a_SN | Zero_b_SN) | Inf_a_SN) | Inf_b_SN) | NaN_a_SN) | NaN_b_SN : ((Zero_a_SN | Inf_a_SN) | NaN_a_SN) | Sign_a_D)} && (Start_S && Ready_SI);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:250:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:252:8
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:254:13
			Special_case_dly_SBO <= 1'sb0;
		else if (Start_S && Ready_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:258:13
			Special_case_dly_SBO <= Special_case_SBO;
		else if (Special_case_dly_SBO)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:262:10
			Special_case_dly_SBO <= 1'b1;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:266:13
			Special_case_dly_SBO <= 1'sb0;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:274:4
	reg Sign_z_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:275:4
	reg Sign_z_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:277:4
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:279:8
		if (Div_start_SI && Ready_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:280:12
			Sign_z_DN = Sign_a_D ^ Sign_b_D;
		else if (Sqrt_start_SI && Ready_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:282:12
			Sign_z_DN = Sign_a_D;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:284:12
			Sign_z_DN = Sign_z_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:287:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:289:8
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:291:13
			Sign_z_DP <= 1'sb0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:295:13
			Sign_z_DP <= Sign_z_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:299:4
	reg [2:0] RM_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:300:4
	reg [2:0] RM_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:302:4
	always @(*)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:304:8
		if (Start_S && Ready_SI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:305:12
			RM_DN = RM_SI;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:307:12
			RM_DN = RM_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:310:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:312:8
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:314:13
			RM_DP <= 1'sb0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:318:13
			RM_DP <= RM_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:321:4
	assign RM_dly_SO = RM_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:323:4
	wire [5:0] Mant_leadingOne_a;
	wire [5:0] Mant_leadingOne_b;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:324:4
	wire Mant_zero_S_a;
	wire Mant_zero_S_b;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:326:3
	lzc #(
		.WIDTH(53),
		.MODE(1)
	) LOD_Ua(
		.in_i(Mant_a_D),
		.cnt_o(Mant_leadingOne_a),
		.empty_o(Mant_zero_S_a)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:335:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_norm_DN;
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_norm_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:337:4
	assign Mant_a_norm_DN = (Start_S && Ready_SI ? Mant_a_D << Mant_leadingOne_a : Mant_a_norm_DP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:339:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:341:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:343:13
			Mant_a_norm_DP <= 1'sb0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:347:13
			Mant_a_norm_DP <= Mant_a_norm_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:351:4
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_norm_DN;
	reg [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_norm_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:352:4
	assign Exp_a_norm_DN = (Start_S && Ready_SI ? (Exp_a_D - Mant_leadingOne_a) + |Mant_leadingOne_a : Exp_a_norm_DP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:354:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:356:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:358:13
			Exp_a_norm_DP <= 1'sb0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:362:13
			Exp_a_norm_DP <= Exp_a_norm_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:366:3
	lzc #(
		.WIDTH(53),
		.MODE(1)
	) LOD_Ub(
		.in_i(Mant_b_D),
		.cnt_o(Mant_leadingOne_b),
		.empty_o(Mant_zero_S_b)
	);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:376:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_norm_DN;
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_norm_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:378:4
	assign Mant_b_norm_DN = (Start_S && Ready_SI ? Mant_b_D << Mant_leadingOne_b : Mant_b_norm_DP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:380:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:382:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:384:13
			Mant_b_norm_DP <= 1'sb0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:388:13
			Mant_b_norm_DP <= Mant_b_norm_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:392:4
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_norm_DN;
	reg [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_norm_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:393:4
	assign Exp_b_norm_DN = (Start_S && Ready_SI ? (Exp_b_D - Mant_leadingOne_b) + |Mant_leadingOne_b : Exp_b_norm_DP);
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:395:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:397:9
		if (~Rst_RBI)
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:399:13
			Exp_b_norm_DP <= 1'sb0;
		else
			// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:403:13
			Exp_b_norm_DP <= Exp_b_norm_DN;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:411:4
	assign Start_SO = Start_S;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:412:4
	assign Exp_a_DO_norm = Exp_a_norm_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:413:4
	assign Exp_b_DO_norm = Exp_b_norm_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:414:4
	assign Mant_a_DO_norm = Mant_a_norm_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:415:4
	assign Mant_b_DO_norm = Mant_b_norm_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:416:4
	assign Sign_z_DO = Sign_z_DP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:417:4
	assign Inf_a_SO = Inf_a_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:418:4
	assign Inf_b_SO = Inf_b_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:419:4
	assign Zero_a_SO = Zero_a_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:420:4
	assign Zero_b_SO = Zero_b_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:421:4
	assign NaN_a_SO = NaN_a_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:422:4
	assign NaN_b_SO = NaN_b_SP;
	// Trace: /vortex/third_party/cvfpu/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:423:4
	assign SNaN_SO = SNaN_SP;
endmodule